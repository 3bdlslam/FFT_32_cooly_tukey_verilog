`timescale 1ns / 1ps


module test_FFT_32;
// Inputs
reg [255:0] Xn_vect_real;
reg [255:0] Xn_vect_imag;
reg clk;
// Outputs
wire [255:0] Xk_vect_real;
wire [255:0] Xk_vect_imag;
// Instantiate the Unit Under Test (UUT)
FFT_32 uut (
.Xn_vect_real(Xn_vect_real),
.Xn_vect_imag(Xn_vect_imag),
.Xk_vect_real(Xk_vect_real),
.Xk_vect_imag(Xk_vect_imag),
.clk(clk)
);

initial begin

/*[(-0.5625-0.5625j), (0.1875+0.375j), (-0.875-0.8125j), (0.4375+0.1875j), (0.8125-0.5j), (0.0625+0.9375j), (1+0.4375j), (0.625+0.1875j), (0.9375+0.5625j), (0.375+0.375j), (-0.5-0.1875j), (0.8125-0.9375j), (0.9375+0.875j), (-0.1875-0.125j), (-0.0625-0.6875j), (1+0.125j), (-0.1875-0.3125j), (0.8125+0.3125j), (0.1875-0.0625j), -0.5625j, (-1+0.5625j), (0.5625-0.0625j), (0.8125+0.875j), (-0.9375-0.625j), (-0.875-0.6875j), (-0.75+0.625j), (0.625+0.125j), (0.75-0.9375j), (0.5625-0.875j), (-0.9375+0.6875j), (-0.8125+0.125j), (-0.4375-0.4375j)]*/
#10 clk<=0;
Xn_vect_real = 256'hF703F2070D01100A0F06F80D0FFDFF10FD0D0300F0090DF1F2F40A0C09F1F3F9;
Xn_vect_imag = 256'hF706F303F80F07030906FDF10EFEF502FB05FFF709FF0EF6F50A02F1F20B02F9;
#10 clk<=1;
/*[-0.8125j, (0.75-0.375j), (-1-0.875j), (-0.4375+0.8125j), (-1-0.6875j), (0.375-0.6875j), (0.6875+0.625j), (-0.5625-0.25j), (0.9375-0.4375j), (1-0.75j), (0.625-0.6875j), (0.0625-0.8125j), (0.3125+0.125j), (-0.125-0.9375j), (0.125+0.5j), (-0.3125+0.75j), (-0.375-0.625j), (0.25+0.75j), (0.8125-0.1875j), (0.8125+0.875j), (-0.625-0.75j), 0.0625j, (0.125+0.6875j), (0.375+0.5625j), (-0.8125-0.4375j), (-0.75+0.9375j), (-0.4375-0.875j), (-0.8125+0.625j), (0.125+1j), (0.9375+0.75j), (0.875-0.6875j), (-0.625+0.25j)]*/
#10 clk<=0;
Xn_vect_real = 256'h000CF0F9F0060BF70F100A0105FE02FBFA040D0DF6000206F3F4F9F3020F0EF6;
Xn_vect_imag = 256'hF3FAF20DF5F50AFCF9F4F5F302F1080CF60CFD0EF4010B09F90FF20A100CF504;
#10 clk<=1;
/*[(0.25+1j), (0.1875-0.625j), (-0.25-0.875j), (0.375+0.5j), (-0.5-0.0625j), (-1-0.125j), (-0.75+0.1875j), (-0.6875+0.0625j), (0.125+1j), (0.5-0.0625j), (-0.25-0.9375j), (0.6875-0.25j), (-0.5625+0.625j), (-0.5-0.6875j), (0.625-0.25j), 0.125j, (0.875+0.0625j), (1-0.8125j), (0.125-0.8125j), (0.125+0.4375j), (-0.625-0.0625j), (-1+0.5625j), (0.875-0.9375j), (-0.5+0j), (0.4375+0.0625j), (0.8125+1j), 0.1875j, (0.5625-0.8125j), (-0.5625-1j), (0.4375+1j), (-0.875+0.5625j), (0.875+0.125j)]*/
#10 clk<=0;
Xn_vect_real = 256'h0403FC06F8F0F4F50208FC0BF7F80A000E100202F6F00EF8070D0009F707F20E;
Xn_vect_imag = 256'h10F6F208FFFE030110FFF1FC0AF5FC0201F3F307FF09F100011003F3F0100902;
#10 clk<=1;
/*[(0.25-0.125j), (-0.625-0.875j), (-0.3125-0.9375j), (0.9375-0.875j), (-1+0.125j), (-0.125+0.5j), (-0.25-0.1875j), (0.625+0.875j), (0.5-0.8125j), (0.1875-0.25j), (0.8125+0.0625j), (0.1875+0.8125j), (-1+0.125j), (-0.875-0.0625j), (-0.75+0.375j), (-0.125-0.625j), (-1-0.1875j), (-1-0.625j), (0.25-0.625j), (-0.0625+0.8125j), (0.25+0.75j), (-0.125-0.125j), (0.5-0.375j), (0.75-0.9375j), (0.375-0.0625j), (-0.625+0.375j), (0.125-0.5625j), (0.875-0.3125j), (0.9375+0.3125j), (-0.0625-0.1875j), (-0.9375-0.3125j), (0.25-1j)]*/
#10 clk<=0;
Xn_vect_real = 256'h04F6FB0FF0FEFC0A08030D03F0F2F4FEF0F004FF04FE080C06F6020E0FFFF104;
Xn_vect_imag = 256'hFEF2F1F20208FD0EF3FC010D02FF06F6FDF6F60D0CFEFAF1FF06F7FB05FDFBF0;
#10 clk<=1;
/*[(-1-1j), (-0.5-0.9375j), (0.4375+0.9375j), (0.0625+0.1875j), (0.625-0.0625j), (0.125-0.375j), (0.875-0.875j), (0.375-0.3125j), (-0.625-0.0625j), (0.1875+0.75j), (-0.625-0.1875j), (-0.25+0.3125j), (0.5625-0.625j), (-0.9375+0.125j), (-0.9375+0.0625j), -0.5625j, (0.9375+0.125j), (-0.25-0.25j), (1+0.125j), (-0.375-0.125j), (0.75+0.6875j), (-0.375+0.875j), -0.6875j, (-0.375+0j), (0.875-0.5625j), (-0.6875+0j), (0.4375-0.5j), (-0.75-1j), (-0.4375-0.9375j), (0.4375-0.6875j), (-0.8125-0.625j), (-0.8125-0.6875j)]*/
#10 clk<=0;
Xn_vect_real = 256'hF0F807010A020E06F603F6FC09F1F1000FFC10FA0CFA00FA0EF507F4F907F3F3;
Xn_vect_imag = 256'hF0F10F03FFFAF2FBFF0CFD05F60201F702FC02FE0B0EF500F700F8F0F1F5F6F5;
#10 clk<=1;
/*[(-0.8125+0.9375j), (-0.4375+0.3125j), (-0.5625+0.5j), (0.875-0.75j), (-0.1875+0.875j), (-0.625+0.375j), (-0.75-0.9375j), (0.9375+0j), (0.6875+0.375j), (-0.125-0.125j), (0.6875-0.75j), (0.5625-0.0625j), (-0.6875-0.75j), (-0.3125-0.875j), (0.4375-0.125j), (0.125+0.125j), (0.625-0.875j), (-0.875+0.8125j), (0.8125-1j), (0.375+0.0625j), (0.0625+0.8125j), (0.6875+0.1875j), (0.8125+0.4375j), (0.8125-0.625j), (-0.9375+0.375j), (0.375+0.125j), (1+0.6875j), (-0.9375+0.1875j), (-0.75+0.25j), (-0.5+0.125j), (-1-0.5j), (0.3125-0.8125j)]*/
#10 clk<=0;
Xn_vect_real = 256'hF3F9F70EFDF6F40F0BFE0B09F5FB07020AF20D06010B0D0DF10610F1F4F8F005;
Xn_vect_imag = 256'h0F0508F40E06F10006FEF4FFF4F2FE02F20DF0010D0307F606020B030402F8F3;
#10 clk<=1;
/*[(0.0625+0.25j), (-0.75-0.6875j), (-0.125-0.4375j), (0.5+0.9375j), (-0.625+0.0625j), (0.6875-0.1875j), (0.4375-0.6875j), (0.625+1j), (0.5-0.3125j), (0.5625-0.875j), (0.0625+0.125j), (0.75-0.25j), (0.3125+0.375j), (-0.0625-1j), (-0.6875+0.5j), (0.125+0.4375j), (0.5625+0.25j), (0.125+0.125j), (0.8125+0.375j), (0.75-0.75j), (-0.875+0.25j), (0.6875+0.1875j), (-0.5-0.9375j), (0.75-0.125j), (0.9375+0.5j), (0.8125+0.6875j), (-0.9375+0.9375j), (0.1875-1j), (0.625+0.1875j), (-0.5625+0.125j), (0.0625-0.3125j), -0.875j]*/
#10 clk<=0;
Xn_vect_real = 256'h01F4FE08F60B070A0809010C05FFF50209020D0CF20BF80C0F0DF1030AF70100;
Xn_vect_imag = 256'h04F5F90F01FDF510FBF202FC06F00807040206F40403F1FE080B0FF00302FBF2;
#10 clk<=1;
/*[(0.9375-0.625j), (0.5+1j), (-0.75+0.1875j), (-0.4375-0.8125j), (0.875+0.8125j), (0.4375-0.5625j), (-0.5625-0.9375j), (-0.125+0.8125j), (-0.3125+0.25j), (0.5625+0.75j), (0.6875+0.0625j), (0.4375-1j), (-0.875+0.4375j), (-0.75+0.6875j), (0.0625+0.8125j), (-0.8125-0.3125j), (-0.375+0j), (-0.1875-0.25j), (-0.4375+0.5j), (0.6875+0.0625j), (-0.5625-0.1875j), (0.25+0.6875j), (-0.9375-0.5j), (-0.5625-0.5625j), (-0.75+0.125j), (0.75-0.125j), (0.4375-0.1875j), (-0.625-0.5j), (1+0.875j), (0.6875+0.4375j), (-0.625-0.3125j), (0.875-0.5625j)]*/
#10 clk<=0;
Xn_vect_real = 256'h0F08F4F90E07F7FEFB090B07F2F401F3FAFDF90BF704F1F7F40C07F6100BF60E;
Xn_vect_imag = 256'hF61003F30DF7F10D040C01F0070B0DFB00FC0801FD0BF8F702FEFDF80E07FBF7;
#10 clk<=1;
/*[(0.375+0.75j), (-1+0.4375j), (0.875-0.625j), (0.25+0.25j), (0.4375+0.3125j), (0.3125+0.75j), (0.9375-0.375j), (0.5-0.3125j), (-0.75+0.5625j), (0.1875-0.4375j), (0.375+0j), (-0.5+0.0625j), (0.9375-0.75j), (0.8125-0.4375j), (-0.125+0.875j), (-0.6875+0.375j), (-0.625+0.5625j), (0.125+0.3125j), (0.0625-0.875j), (0.125+0j), (0.875+0.125j), (0.8125+0.1875j), (-0.25+0j), (1-0.625j), (1+0.5j), (0.25-1j), (-0.4375+0.25j), (0.25-0.5625j), (0.8125+0.875j), (-0.8125-1j), (-0.4375-1j), (0.5+0.75j)]*/
#10 clk<=0;
Xn_vect_real = 256'h06F00E0407050F08F40306F80F0DFEF5F60201020E0DFC101004F9040DF3F908;
Xn_vect_imag = 256'h0C07F604050CFAFB09F90001F4F90E060905F200020300F608F004F70EF0F00C;
#10 clk<=1;
/*[(0.25+0.0625j), (-0.9375+0.625j), (0.125+0.3125j), (0.8125-0.1875j), (-0.375-0.3125j), (0.0625-0.625j), (-0.25+0.8125j), (-0.125-0.375j), (0.375-0.625j), (0.8125+0.875j), (0.125-0.75j), (-1+0.3125j), (0.9375+0.375j), (-0.25+0.8125j), (0.875-0.8125j), (-0.875-1j), (0.875+0.9375j), (0.125+0.6875j), (0.6875+0.0625j), (0.5+0.625j), (0.625-0.6875j), (0.4375-0.25j), (0.375+0.625j), (0.75+0.0625j), (0.625-0.3125j), (0.1875-0.625j), (-0.625+0.25j), (-0.75+1j), (-0.5-0.375j), (-0.25-0.6875j), (0.4375-0.1875j), (0.125-0.3125j)]*/
#10 clk<=0;
Xn_vect_real = 256'h04F1020DFA01FCFE060D02F00FFC0EF20E020B080A07060C0A03F6F4F8FC0702;
Xn_vect_imag = 256'h010A05FDFBF60DFAF60EF405060DF3F00F0B010AF5FC0A01FBF60410FAF5FDFB;
#10 clk<=1;
end

always @(Xn_vect_real,Xn_vect_imag)
$monitor("input:\nreal=%h  imag=%h\noutput:\nreal=%h  imag=%h",Xn_vect_real,Xn_vect_imag,Xk_vect_real,Xk_vect_imag);


//Expected output:
/*[ 3.375     -1.j         -1.12500074-6.12111192j  0.01204895-2.77623195j
 -6.55007451+0.48599221j -5.01332521-0.35799513j -0.62408572-2.29758482j
  4.77055505-3.25459845j -1.22802651+1.8779878j   6.375     +1.375j
  7.07705696-4.45957884j -3.64142962+5.10977216j  1.33196161-0.1625996j
 -0.75444174-5.83286886j -0.01862674+4.67797528j -3.57258112-4.06199985j
  3.00415273-4.51723568j -1.375     -1.25j        0.95398024-3.08369053j
 -4.95919451-1.80111743j -3.88609526+3.66158985j -2.36167479+1.23299513j
  0.86819472+4.8247406j  -0.06820567-0.47135303j -1.19849905+2.31476591j
 -5.875     -2.875j       2.60437118-8.72775432j  5.58857517+3.21757722j
  0.48288782+4.03278449j  0.12944174+0.70786886j -2.73588991-1.31299543j
 -4.62976826-1.96204867j -4.95630683+4.80671502j]*/
//real=36EE0098B0F74CED6671C615F400C730EA0FB1C2DB0DFFEDA229590702D5B6B1  imag=F09FD407FBDCCC1E16B951FEA34AC0B8ECCFE43A134DF925D28033400BEBE14C
//real=36ecfd9bb0f348ed666bca13f400c72aea12b5c1da1300eba22b540502d6b9ba  imag=f09fd207fadecd1f16b84f01a444c0bfeccde6371446f523d27c353d0af0e24b

/*[ 1.3125     -1.5625j     -7.60248489 -3.89058697j
 -0.04619098 +1.67479848j  2.43194221 +2.95470782j
 -2.19378157 +0.07766504j -0.4425499  -0.3418908j
  1.15368711 -4.44449351j  4.5069385  -1.36189146j
 -6.3125     -5.0625j     -1.97751231 -0.5426202j
 -3.91261647 +2.48825819j  1.66829908 +0.71450489j
  6.27849026 -5.22671356j -1.59915321 -1.13191353j
  1.05449616 -6.6323967j  -5.51890235 -0.23443734j
 -0.5625     -6.6875j      4.67566712 -3.09066863j
 -3.51554693 +0.70648308j -1.09660968 +4.11511266j
 -3.43121843 -0.45266504j  3.85462498 +1.82762741j
  6.06490505 +1.4042022j  -0.44380436 +8.16208571j
 -0.1875     +2.8125j      2.51524279 +2.95585631j
 -4.77564561 +1.13046024j -2.21073838 -3.65564571j
  3.09650974 -2.39828644j  3.57616542-11.28580359j
 -0.02308833 -0.82731199j  3.66287499 +1.80556343j]*/
//real=15870026DDF912489BE1C21A64E710A8F74AC8EFCA3D61F9FD28B4DD3139003A  imag=E7C21A2F01FBB9EBAFF8270BADEE96FD95CF0B41F91D167F2D2F12C6DA80F31C


/*[ 0.8125    -0.8125j     -1.9907069 +5.12987704j  2.44858062+1.75142617j
 -1.56650586-0.27580098j  2.51202426-2.38410669j -3.93063964+3.53920576j
 -4.46123826-2.01881112j  0.0870567 -2.84979285j  0.        +5.5j
  6.67800648+1.15169779j -0.42149554+3.82708393j  0.21007052+8.09254971j
  2.97649035-1.73505817j -0.11971167+3.20885238j  0.28810141+5.06544303j
 -7.50132644-0.24982255j -2.9375    -1.6875j     -0.09604306+0.60665449j
 -4.00556114-2.28175625j  0.05164287-3.45010324j  1.36297574+8.13410669j
 -0.64162912+1.5053089j   2.61136452+1.13492764j -1.48614537+1.47408828j
 -0.125     +3.5j         1.60849094-6.83797679j  5.22847606-3.29675384j
 -0.70256683+2.3759952j   8.89850965+6.48505817j  0.99223296+1.69638043j
  2.81177233-4.18155956j -1.59222558-0.11711357j]*/
//real=0DE127E728C2B901006AFA032FFF0488D1FFC00015F629E9FE1953F57F0F2CE7  imag=F3521CFCDA38E0D358123D7FE53351FDE509DCC97F1812173893CC26671BBEFF


/*[-1.0625    -4.9375j      4.28050011-1.137117j   -7.01084847-3.60743189j
  0.02349401+2.58679867j -1.11113591-7.06640287j -3.6810547 +0.56075969j
 -1.38467298-0.46765064j  7.9906515 -2.33258944j -0.125     +9.375j
  2.29234966+5.36543744j  2.12560495+2.47856757j  0.61159533-2.04571669j
  3.87001939+2.6851213j  -0.63162297-0.75632708j -0.32575436+3.1419985j
  0.25786183-1.95285639j -1.4375    +0.0625j     -4.15499416+3.12109474j
 -1.90488926+4.16288824j  4.00836323+3.60282744j -0.13886409-2.55859713j
  2.84675196-3.97280049j -0.97256006-0.48945614j  2.40501983+0.16616986j
 -0.125     -4.j         -0.771409  +0.17875941j  2.04013277+1.96597608j
 -0.88609326+6.8591389j   1.12998061-3.0601213j   3.8194791 -3.85980671j
 -5.5670126 -2.68489171j  1.58910753-5.38377236j]*/
//real=EF449000EFC6EA7FFE2422093DF6FB04E9BEE240FE2DF126FEF420F2123DA719  imag=B1EEC7298F08F9DB7F5527E02AF432E101314239D8C1F902C0021F6DD0C3D6AA


/*[-2.0625    -6.875j      -0.07868576-5.49224583j  2.17587352-6.41779889j
 -3.29911183+2.86932925j  1.58524756-2.90847087j  0.42441627+0.24747381j
 -3.69085483-4.9221665j  -5.20075794-4.78442871j  3.        -0.8125j
 -4.01518385-1.95594554j  1.24508188+0.21124617j  1.07353089-2.42806395j
 -3.41475244+3.19768443j -2.02117835+0.92887454j -1.63139065+7.6440932j
 -2.72012355-2.44034344j  6.1875    -1.5j        -2.95249904+4.22313805j
  1.22057309+1.29647855j -1.8425298 -5.70778575j  0.78975244-2.46652913j
  5.50114135+3.34984264j  1.16572856-2.97732843j  0.05800259+0.29362176j
 -0.375     -0.5625j     -3.12304873-0.75502424j  2.85847151-1.08992582j
 -3.73734561-4.70314947j -4.21024756-0.07268443j -5.23496189+2.45388656j
 -5.84348309+4.25540173j -3.83166474-4.0991797j ]*/
//real=DFFF22CC1906C5AD30C01311CAE0E6D563D113E30C581200FACF2DC5BDADA3C3  imag=92A99A2DD203B2B4F3E103DA330E7AD9E84314A5D935D104F7F4EFB5FF2744BF


/*[ 6.87500000e-01-0.625j      -8.45260488e+00+2.78397661j
 -8.82143345e-01-3.86883157j  2.01900619e+00-0.89231345j
  3.85301452e+00-1.26570392j  2.46792013e+00-1.96383122j
 -1.77492242e+00+5.15479544j -9.74605645e-01+3.97137248j
 -6.25000000e-01+8.5625j      7.46769530e+00-0.67211345j
  6.62826835e+00-3.35894338j -4.49847359e+00+3.44116468j
  1.31380096e+00+2.81380096j -8.01217112e+00+1.43713836j
 -7.69194432e-02-2.72971951j -2.22945061e+00+4.0325233j
 -1.81250000e+00+1.25j       -6.10545252e+00+4.90206754j
  2.02338613e+00+0.22238496j -3.64259318e-03+5.72488155j
 -4.78014517e-01-4.35929608j  1.88488485e+00-1.72503633j
 -2.03844165e-04-1.96025179j  1.37526057e+00+5.43121283j
 -6.25000000e+00-1.1875j     -2.19517180e+00-2.72839679j
  1.23048886e+00-0.99461001j -5.03465697e+00+3.00139348j
 -1.88800955e-01+1.31119904j  1.44490004e+00-0.53380472j
 -6.64795429e+00+2.03517586j -2.15343736e+00+2.78976512j]*/
//real=0B80F2203D27E4F1F6776AB91580FFDDE39F2000F91E00169CDD13B0FD1796DE  imag=F62CC3F2ECE1523F7FF6CB372D16D540144E035BBBE5E156EDD5F13014F8202C


/*[ 5.8125    -1.125j      -3.23132829-1.96126597j -3.58566902-1.45971212j
  1.17949843-2.38646158j  3.60409226-0.02458739j -1.39214668+3.97336212j
 -3.05022577-3.70133326j  0.33537983-5.78697716j  1.375     +4.1875j
  0.48716923+8.56163173j -0.02662454+6.50979161j -0.54609379+2.4336535j
 -0.29863591-1.32268443j -0.47020758-0.79028961j  8.36535686-0.64193374j
  3.21805509-0.94343429j -4.5625    +3.375j      -0.03183131-2.08355856j
 -1.27936975+4.92678013j -0.94749604+3.52420657j  6.52090774-1.35041261j
 -1.56980824+5.1515365j  -3.64324013-4.52614238j  0.44004108+4.19418831j
  3.375     -0.1875j     -0.88301937-3.65069068j  0.64166332+1.02314038j
 -0.02689885-4.08396163j  0.67363591+1.94768443j -3.40882776-5.70072553j
 -3.92189096+0.36940939j -1.15248574-0.45121372j]*/
//real=5DCDC71239EAD005160700F8FCF97F33B700ECF168E7C60736F20A000ACAC2EE  imag=EEE1E9DA003FC5A4437F6826EBF4F6F136DF4E38EB52B843FDC610BF1FA505F9


/*[-5.00000000e-01+1.0625j      6.36130349e+00-1.98832231j
 -9.33441001e-01+2.37354622j  7.34279144e-05+3.62476237j
 -2.77189303e-01-4.14330583j  5.47166347e+00+1.7661857j
  3.93283846e+00-0.38719347j  3.67463303e+00-0.69958635j
  7.56250000e+00-0.75j        6.54632819e+00+1.0737701j
  3.76274573e+00-1.35944232j  1.64845131e+00-0.38228198j
 -3.71913104e+00-2.61817956j -7.03969288e+00-0.67190084j
  2.73366617e+00-1.3392808j   5.90389023e-01+0.25732234j
 -3.87500000e+00+1.5625j      5.17091611e-01-2.10923263j
 -7.27092905e-01+3.73673515j -8.65686945e-01-5.4584118j
  1.40218930e+00-4.23169417j -5.43559375e+00-6.92751098j
  1.04571493e+00-0.53069975j  4.61694823e+00+3.4792813j
 -3.43750000e+00+4.875j       3.28543181e+00+4.07708569j
  1.64778818e+00-9.50083906j -3.81101239e+00-1.36249571j
 -1.15586896e+00+2.24317956j  1.79346806e+00-3.72007474j
  1.53778044e+00-0.99282598j  3.64620431e+00-0.95859017j]*/
//real=F865F200FC573E3A79683C1AC5902B09C208F5F316AA1049C9341AC4EE1C183A  imag=11E12539BE1CFAF5F411EBFAD7F6EB0419DF3BA9BD92F8374E4180EB23C5F1F1


/*[ 6.1875     -0.0625j      1.6053308  +0.82967418j
 -1.8065116  -0.41981846j  2.87068693 -3.38209808j
 -4.51960678 +3.18382034j  5.29723842 +1.69938816j
 -3.81644818 +2.73311992j  2.23732966 +3.54127451j
  0.9375     +5.4375j     -3.10717642+11.11099145j
  1.0092     +0.53468278j -3.64734725 -1.53911482j
 -2.4892767  +4.33026695j -0.06115936 -1.12982894j
  6.32287615 -4.72209282j  5.30643722 +1.15016296j
  1.9375     +2.4375j     -0.62631065 -1.60430555j
 -1.75046891 -3.5084824j   1.86149229 -3.42496876j
 -3.10539322 -1.05882034j  4.37125722 -0.36483592j
 -0.28342555 -4.1687801j   0.13577027 -6.00323068j
  3.1875     +3.9375j      0.72130202 +3.42404757j
  1.79778051 +6.14361808j  0.19029429 -2.14645903j
 -2.1357233  +0.79473305j  0.29951796 +1.53486906j
 -5.47300241 +5.40775299j -1.45466341 -0.6955661j ]*/
//real=6319E42DB854C3230FCF10C6D90065541FF6E41DCF45FC02330B1C03DE04A9E9  imag=FF0DFACA321B2B38577F08E845EEB51227E7C8CAF0FBBEA03F3662DE0C1856F5


/*[  4.1875    +0.3125j      -3.97906721-0.52487417j
   0.13648719-2.54850139j   3.06860751+0.72603631j
   5.25022321+1.52458739j  -1.40250694+3.12023639j
   1.19725225+4.63374751j  -3.19902285+3.73666955j
   1.75      -2.j          -2.80758653-3.38033655j
   0.76327978+5.36865866j   4.11015089-0.4557042j
   5.66811643+0.7771893j   -0.76237555-1.9633596j
   1.76306763-2.9578805j   -2.82964747+2.75745225j
   4.9375    -1.5625j      -4.44054341+0.51618895j
   6.33362914+4.41201601j   3.04878109-4.2623018j
  -3.50022321+2.85041261j  -0.46268868-1.37002924j
   2.20179626+0.89918449j  -1.35229128-8.55924257j
   0.375     -0.5j          3.76488654-1.40907527j
 -10.73339611+1.26782673j  -1.40126785-0.684807j
  -1.66811643-0.9021893j    2.58988177+0.0112495j
  -0.66211615+4.4249485j   -3.94531003-2.25810255j]*/
//real=43C1023154EA13CD1CD40C415AF41CD34FB96530C8F923EB063C80EAE629F6C1  imag=05F8D80B18314A3BE0CA55F90CE1D12CE70846BC2DEB0E80F8EA14F6F20046DC


endmodule