`timescale 1ns / 1ps


module test_FFT_32;
// Inputs
reg [255:0] Xn_vect_real;
reg [255:0] Xn_vect_imag;
reg clk;
// Outputs
wire [255:0] Xk_vect_real;
wire [255:0] Xk_vect_imag;
// Instantiate the Unit Under Test (UUT)
FFT_32 uut (
.Xn_vect_real(Xn_vect_real),
.Xn_vect_imag(Xn_vect_imag),
.Xk_vect_real(Xk_vect_real),
.Xk_vect_imag(Xk_vect_imag),
.clk(clk)
);

initial begin

Xn_vect_real = 0'h03F5F1020B02F60DF005090D04F60DF4FDFD0FF4F80306FD010FF0F8F6F0F301;
Xn_vect_imag = 0'h0A0F08F4F5F90DFBF00E07F3F30C05FD080B0A0B060FFF0D0EFA050009F204F9;
#100;

Xn_vect_real = 0'h0C05FB060A10070F04F0F1F20DF2030608100C0CFC0010FFFB020608FDF4F2F4;
Xn_vect_imag = 0'h0EF80801FEF70A0600FD0003F910030DF9F11006FCFE0EF5000D08FD10F7F203;
#100;

Xn_vect_real = 0'h070F00FBF2FC0801FEF1F1090FF1FFFF040B0500FA02F1FBFAF7FEFCFC0DF3F8;
Xn_vect_imag = 0'h0EF3F20EF1F710F7F3F10F0200FDF809F609000FF3FC02FD10F8040CFE0208F3;
#100;

Xn_vect_real = 0'h08F3100D030CF4F104F40E0C070FF204F9FE0E05F2F8F60FFF02010CF208F308;
Xn_vect_imag = 0'h10F2F3F9F101000AFF0710F6F4F8010F08FA01FEFEFBF6FCF7F904020D0CF4F7;
#100;

Xn_vect_real = 0'h080910F910FBFA100AFF05FBF90AF005F4F7F2F1F1F70000F108FB0E0909FF00;
Xn_vect_imag = 0'hFD080308F805F60AF50F0F0C0FF908071002F20A0A060E0AFF04FF08100D1009;
#100;

Xn_vect_real = 0'hF4F6FDF2FC0E090D0BF8FBFE0DF302020E0AFB0C030A00F2F70BF108FDF9F1FF;
Xn_vect_imag = 0'h0106FB0406FD00FEF0F1FDFBF80F01FE10FEF810100AF5F3F504F0F3FAFFF6F2;
#100;

Xn_vect_real = 0'h08FC0300FEF7FBFCFAF1011003F2F200F30CF70B0B03090E0DFF020208100702;
Xn_vect_imag = 0'h070C05F4FA0EFD07FB0802F604F609F608F902030B0DF9F00BFF0902FD05F1FA;
#100;

Xn_vect_real = 0'h0600F8FBF0FAF505FB0D090E0D0FF00AF005F00FFB0FFBF507F0F0F50AF40AFD;
Xn_vect_imag = 0'h0B010B0A0CF1F80710F00B070206F503F50AF40B0C100E0608FE04F7F707F1F7;
#100;

Xn_vect_real = 0'h0B03F20006FFF6FF0403F9FEFA04F2070B050507F70EFDF00DF4F80003FAF0F0;
Xn_vect_imag = 0'h02FFF506080C05FBFF0906FB04FA0D04F2F7FFF6050EF0F8F1040DFE040FFAFF;
#100;

Xn_vect_real = 0'hFAF7F010FDF50F10F4FBF1FF09F70FFBF1F8F6F4F20A0F02F1F305F8FE0E09F1;
Xn_vect_imag = 0'hF210FEFCFCFEF30AFB01F30E090FFDFDF203F10F0204F0FD05FB0E00FE0C030F;
#100;

end

always @(Xn_vect_real,Xk_vect_imag)
$monitor("real=%h  imag=%h",Xk_vect_real,Xk_vect_imag);


//Expected output:
//real=CE88FA161E1F3C5731250319E10C77D5F8AF3E05DCB2E17FC1E5FDDEF622AB0D  imag=52A801F228662957DDE71EEBEAE6162C224C14B10F0D08AFCB21F8CD42412BFD
//real=3EDC05B816643D1EF61AABFEDE5ACE101CC7351E160E6C2A3C113205028419EC  imag=38FC87E0003CB850F4123DD3EB13C93A36212DDE24E6227FC6F2394D010869ED
//real=CAC925EE1AF03BF1D7F2E87F3EF423DBE8F2CDE0E407F5445FA20A67F4FA6023  imag=F2E6FF00DC07ADE1C7F0303A5362A45F0E1AD0245C343643DD347FFD08DC0100
//real=2617D9BCD72BDB70E7E6F61510351111B6FDE22D7F0C0BFC05EC00BEE26448FF  imag=D8D90E87D6391F473F1B5F417F09423F0AC1F342AB082F37D70D379D7209E803
//real=F963AFE4FFFEF734F31A0DADFE094851D117CD51B8C613162BE207DC1C0B267F  imag=7FCA382AE580F8EDFFBC09D6080A6500C9AEE328AAEF2DFB07C344F6EA40D62B
//real=F8BA2DD0EF44180158E5FCD60E3C09CBE2F21113EFC1B4180292541100A69BA9  imag=BBA2232FD918F2D02F0D7FEC001C0149D9BF25C333A8151A35D71233ADC87CE4
//real=2D1411300013F71068110036DAD3F74EF31EB77B2012FB18D09D18ABBF4ED922  imag=1568F70FFA70FED94EF3CF29121A1EC625B81CE524E60D05E4254A090BE9F297
//real=E1BE497F022F14E21C0D2DD1DE04CE4EA97FEA312DFCB7EA420AECDFCB52BCD9  imag=44BB117FF8F5DFB72F6248C913338004027CF923283F03202FE6FDF3E929A816
//real=D3F1F8DC0211C92E7F39FAF429F7090BE945C8F06DEC012129146FCE1AF82CA9  imag=0D1FC6F399F70815D7291408EBFBFEBBEB060FE1E07FF23D150C2627DAD71828
//real=B20C9FF4C8E6F9CDB45E6851E1B0281DFECBFB2A065F0131B4D5F3EABAFB1821  imag=1404171C482BA1FF2EBFD6D1B1EA9600801DFEAB291FF7FAFEA60466802E0421
endmodule