`timescale 1ns / 1ps

module Test_FFT;

// Inputs
reg [511:0] Xn_vect_real;
reg [511:0] Xn_vect_imag;
reg clk1,clk2,rst;
// Outputs
wire [511:0] Xk_vect_real;
wire [511:0] Xk_vect_imag;

// Instantiate the Unit Under Test (UUT)
FFT uut (
.Xn_vect_real(Xn_vect_real),
.Xn_vect_imag(Xn_vect_imag),
.Xk_vect_real(Xk_vect_real),
.Xk_vect_imag(Xk_vect_imag),
.clk1(clk1),.clk2(clk2),.rst(rst)
);

initial begin;
clk1<=0;
clk2<=1;
rst<=0;
#1 rst<=1;
#1 rst<=0;
end

always begin; #0.06172839506172839; clk1<=~clk1;
end
always begin; #5; clk2<=~clk2;
end

initial begin;

#10;
Xn_vect_real=  512'h00AF_0099_00A5_008C_0044_00DA_00FF_0069_0090_0079_00DF_0056_00D0_008E_005E_0028_0010_00F6_00DD_00E8_00ED_0001_0035_000D_0031_0062_0095_0037_0040_0053_00BD_0030;
Xn_vect_imag=  512'h0010_00A4_0004_00E4_00C7_00CE_00CC_0033_00D5_00B2_00C2_003E_008F_0002_00A9_00B1_0047_0029_00E9_0055_0036_001A_0074_0098_00F7_0004_0011_008D_0057_0094_0023_008B;
#10;
Xn_vect_real=  512'h00D8_00CC_0059_00E3_00AC_00AC_0019_0046_0013_0030_00DA_00E5_0053_00F7_0014_0006_0035_00AC_00A9_00A6_0077_0044_00B5_00CA_00F9_00F9_00AC_00BA_0051_0045_0003_0015;
Xn_vect_imag=  512'h0016_005C_00C6_00A3_0090_00C8_00DE_00C8_00A0_0056_001C_0043_00B4_0006_00EE_0037_0064_00BD_008D_005B_000B_006F_0015_0060_005B_000D_00F6_00C2_00E9_004B_0083_00CB;
#10;
Xn_vect_real=  512'h0014_0043_0050_00E8_00D8_00A8_00F0_00F1_00E0_00EC_005F_0001_00A6_00A0_00F6_000F_00B4_006B_006C_0052_00EF_0027_00BC_00D8_003C_00FB_0053_005F_00AC_0065_003D_00B9;
Xn_vect_imag=  512'h00C3_0070_0003_00B4_0018_00E5_004B_0080_0058_001E_0074_00B6_008B_0073_0090_0077_0096_0062_0038_007A_0048_000E_00D9_00DA_004E_0055_00BF_0012_00FC_00BE_0032_001D;
#10;
Xn_vect_real=  512'h0037_00B5_0017_00A0_0007_0035_003C_00E1_00D4_00B7_0098_0099_0010_00AB_002C_00EB_0029_00CE_00D4_00F4_005B_0018_009B_00A0_0001_00C7_00C4_003C_0063_0026_0077_00FE;
Xn_vect_imag=  512'h0086_00C2_00FC_00F0_0002_0027_002A_00D4_001F_00F0_00A8_008D_00A3_000B_0028_0014_00B1_00C3_000F_0015_004D_0011_0006_0042_0000_007B_0006_00F1_00E4_0079_00FD_0088;
#10;
Xn_vect_real=  512'h00A4_0016_00E2_0089_0027_001E_0024_0037_0001_00A0_002C_00D4_002A_006A_00F4_0021_00A6_00B4_0006_00CA_00C5_009D_00F6_0076_004A_0095_001B_0054_00DF_008D_003B_0083;
Xn_vect_imag=  512'h00E8_005E_00EF_0097_00D6_00A4_00AE_0036_0049_00EA_006A_00CE_0067_0066_0035_0008_0068_00B7_00B6_007B_00A8_007D_0025_00B8_00A6_0092_00AF_0019_00B8_0035_0086_00C4;
#10;
Xn_vect_real=  512'h00F3_001B_00D4_001E_001F_00EF_0039_00AB_007D_001C_00B4_0089_00A2_0039_009E_0004_00BF_00EF_00F5_00F4_0003_0028_0098_0014_00EC_00D6_0071_00EB_009A_0023_005F_0050;
Xn_vect_imag=  512'h00D7_0019_00B4_0010_0080_0047_005D_00F1_00A6_00A2_00AE_0006_006A_006A_00A4_0029_0022_00E5_0017_00D1_002A_008B_00D4_0056_0004_00BB_00F7_0003_0001_00A4_005A_0083;
#10;
Xn_vect_real=  512'h0077_0074_00D1_0062_00B6_00C3_00F8_00C4_007E_008B_0076_007C_0006_008D_00D0_0062_0070_0097_006E_0003_00B0_005B_009C_0095_00A0_0088_00D6_0053_006C_00D7_0096_00D8;
Xn_vect_imag=  512'h00A8_0020_0049_0051_00DF_0078_0007_00F7_00A2_00D4_0044_00DF_00E4_00CE_00E6_0001_0098_0028_009D_009E_0036_008C_006D_009A_00CF_00ED_0085_0074_00E2_0016_00B7_0072;
#10;
Xn_vect_real=  512'h0075_0070_0082_00A1_009B_004C_0045_00D2_00F7_006B_00C1_00F8_00EF_00EA_000B_00DB_0088_00D1_0006_005C_007C_004C_00CA_00DF_00A1_0097_007D_0080_009C_006B_0099_003C;
Xn_vect_imag=  512'h00C8_008D_000B_00A0_00FF_00B2_007C_0021_0049_0090_0087_0071_0062_0003_0013_000D_00F1_0006_002C_00A8_00F8_008C_008D_00DD_0050_00FB_0043_0071_00AE_0027_0001_00B2;
#10;
Xn_vect_real=  512'h0059_0064_0018_001D_0096_0042_00B9_006A_00EC_00B5_00EE_00C2_001F_0037_006E_00BA_008E_001B_00A4_0005_0038_00F7_009F_00A8_0051_0090_00F1_00BE_00EE_0030_00FC_0054;
Xn_vect_imag=  512'h007C_007B_002A_00F4_00A7_0057_003B_005E_0064_001E_003A_00DC_0054_0068_0032_0094_0019_005C_00D8_00AA_00A5_00BB_0075_0075_00E3_00E0_00E3_005A_00B2_009C_0048_00CE;
#10;
Xn_vect_real=  512'h007A_0013_00F6_00F3_001A_00EC_0084_0037_008E_00D1_0050_0097_0011_0042_00A9_00E5_007B_00E8_00E9_00F6_0048_00F9_0068_006A_00E0_0051_0075_00D4_00A5_00FF_0041_0053;
Xn_vect_imag=  512'h0097_009F_0003_001C_00A2_00D6_006E_00F2_0076_0031_00F9_0046_0002_00E9_0017_00CF_0001_005A_0061_0015_00E0_0069_0076_00F6_0063_003D_00CD_00DA_00C9_001E_00D1_00F8;
end

always @(posedge clk2)
$monitor("real=%h  imag=%h\n\n",Xk_vect_real,Xk_vect_imag);
endmodule

/*
Expected Output:

real=0FFB01B001E5002FFE970183FF160135FD72FF39FFBE02D9FFEB0255FF25FFF0021100F6FEFE01E0FF50FF6A0191FE6DFF86FED9FFB403C8FF2CFFEFFFD2FDC5  imag=0EDEFE09FD7700E7FE4BFFB7FE7F022AFEE30070FE4001EAFF8EFECBFCE0FCF300C6FD00FEA7008600E700D7FF22FFD901910372FF4CFC930240FD0D0030025F
real=0ffb01ab01e3002cfe960182ff140134fd72ff3bffbe02daffea0254ff23ffed021100f7feff01e2ff50ff6a0192fe6cff86fed7ffb403c8ff2cfff4ffd3fdcb  imag=0edefe08fd7700e7fe4affb6fe7f0228fee3006efe3f01e5ff8dfecbfce0fcf300c6fd02fea5008700e800d4ff21ffd801910370ff4dfc950241fd1300300265

real=106D0128FE930062FF1A012201BB002EFF4A005800F0FE2A0142FF8801F6FFD8FE2D0070FD5802EA018C000501B20210019C0320FF220054FF60017EFEA9FF10  imag=0FA7034EFF6CF9A0FBF302C4FF15FFF7FE6AFFD8FC3B00DEFF13FD46005DFE8A0145007AFF5BFF98FF4200FFFF92FF0EFF5E003200FFFE7202ADFFE500F4004B


real=11DEFF85FCBCFF48FEF3FFA2FFE20194003501440212FD41FD74007A032AFF2900B6FB78FEDEFE9EFDB4020C018DFDDD012BFF71FC69009A0112FD77FEB30056  imag=0E87FE7BFE4BFF77010BFEAC017302720054025A02C0028CFF71FFE6002E0014FFEDFEECFF9001130206FEE6020CFFB700D0FF6E005DFFC9FDDEFFA400F1016B


real=0FBD0025FDD6FED204F101F2009F0054FDC0FE680107FF4A0013FFD3FF5D00C9FBD9FFF4FD10FFE4FC97FEBD00F802C7FED200A4FD5F0034FFE501C00217FD60  imag=0E1B02E901C80295FF0FFDD600BAFF6401D2FD8E007C0090FEB3FF570224FE42FE5900A202BD0373FE58FE8DFFCDFFDFFE6AFCACFFA2FDFC01E7FE9401710328


real=0E7FFF2B029801D700F6FC61FF85FF9D00ACFF530071FE30FFD0FFC20179018AFF850005020DFFEB00A900D301A20243FF78FFE1006100D6FD1101B0FFE0FEA6  imag=1128036A000000A3001CFECA0002000600AB014B00C304A2FD15002001CF011D0128028600D9FC64015BFDC9FF1CFDCF0075010E005A018AFFFC014B0022FF93


real=103DFF9E0092FD6700F4023FFFE5FEDF011B01B8FF80FBF001BDFFA30273FEC3022D015900B705CE0307FF9FFE1EFFCFFE5F02FD01560106013AFF84FFB3FEF4  imag=0E6F00D3FF550126FF1A0332FDE9FFABFE4301A6038300D4FF350349FEC501D4003F01B90157FF96FFC3FE82015300A0FDEFFFC10174FF580427002DFED3FF2A


real=11C9021DFD9EFFAD00BFFF0BFFBFFE01FE030071FFB300A80020FE8A00DD00C300FBFEADFEC50014FED70096000DFFE3FEAD0142004B011900FDFE29013D0178  imag=1183FEF4FDAD002C016F0166FEE9009700F30244FE37FFC900BAFF8404F1FFDC0115016501A7FE07FF1BFC8500A1004602A50112FDE100F4FE140072FE91FFC8


real=121DFDDB00A00141011CFDBEFDF5FF43015DFFA8FFF8FE53006502A2FEBE00C7FF4302EAFEEA008AFE920038012BFFBF021FFDD501AEFF82FFB90056FC1C0037  imag=0EE4FFFD001FFFA7FF6AFFDF00E001FD0448FEF7010AFF5CFF29FDB50190FE3F000AFEC101480002FF07FEC9030C0098022EFFFA03DDFF83FF9401FFFD33020D


real=1082FD93FDD9004D01F3FD35011AFFFDFD840145FE11FF9CFF24FEED0048025D0236000D00ABFD2A0088FFB4FF56006FFFC00099032BFFBEFF85FF0DFCD802B6  imag=106B012A017C01B8FF53FFC30075FFDB014301CEFF95FF4F0041FC61FE450050FE83FF77FEE10134000F0202FFD1037A0087FF00FE4301EBFE85FEADFDB30022


real=1265FE99FFF9FD45FD98FE26FE400062FDAEFF57010C02C1006A0331FFD30213FD85FFA10015FDB405BA017CFBDA0159005400F6FFDFFDF4016FFF370153FFE4  imag=106102B1FD810101FF15005B01F100E0FFB2003F01B8FF3DFE93026FFE890091FF07012BFF25FF9FFD98FE1CFD43FE8CFFDE032B01ED01D40151FF12FFF10070


*/
