`timescale 1ns / 1ps


module test_FFT_32;
// Inputs
reg [255:0] Xn_vect_real;
reg [255:0] Xn_vect_imag;
reg clk;
// Outputs
wire [255:0] Xk_vect_real;
wire [255:0] Xk_vect_imag;
// Instantiate the Unit Under Test (UUT)
FFT_32 uut (
.Xn_vect_real(Xn_vect_real),
.Xn_vect_imag(Xn_vect_imag),
.Xk_vect_real(Xk_vect_real),
.Xk_vect_imag(Xk_vect_imag),
.clk(clk)
);

initial begin

/*[(0.9375-0.625j), (-0.125+0.125j), (-0.25-1j), (0.625-0.25j), (0.625-0.6875j), (0.3125+0.4375j), (0.75-0.3125j), (-0.5625-0.9375j), (-0.125-0.125j), (1-0.1875j), (-1-0.0625j), (-0.25+0.625j), (-0.0625+0.0625j), (-1+0j), (-0.75-0.5625j), (0.25-1j), (-0.125-0.75j), (-0.875-0.25j), (0.625+0.9375j), (0.375+0.0625j), (0.4375+0.875j), (-0.125+0.6875j), (0.3125+0.75j), (0.375+0.0625j), (-0.4375-0.5625j), (-0.75-0.0625j), (-0.25-0.125j), (0.125-0.1875j), (0.375-0.5625j), (-0.3125+0.25j), (0.3125+0.6875j), (-0.5-0.75j)]*/
Xn_vect_real = 256'h0FFEFC0A0A050CF7FE10F0FCFFF0F404FEF20A0607FE0506F9F4FC0206FB05F8;
Xn_vect_imag = 256'hF602F0FCF507FBF1FEFDFF0A0100F7F0F4FC0F010E0B0C01F7FFFEFDF7040BF4;
#100;

/*[(-0.5625+0.3125j), (0.8125+0.4375j), (-0.1875-0.75j), (0.375+1j), (0.625+1j), (-0.25+0.5j), (-0.875+0.9375j), (0.625-0.125j), (-0.75+0.1875j), (-0.0625-0.125j), (0.3125+0.75j), (0.3125+0.6875j), (0.875-1j), (0.4375-0.4375j), (-0.125+0.6875j), (-0.75-0.3125j), (0.125+0.5625j), (0.75-1j), -0.4375j, (-0.5-0.625j), (-0.0625+0.5625j), (-0.1875+0.1875j), (0.4375-0.4375j), (-1+0.0625j), (-0.5625-0.1875j), (0.5+0.5625j), (0.1875+0.0625j), (-0.5-0.5625j), (0.6875-0.1875j), (-0.875+0.3125j), (0.625-0.8125j), (-0.125+0.375j)]*/
Xn_vect_real = 256'hF70DFD060AFCF20AF4FF05050E07FEF4020C00F8FFFD07F0F70803F80BF20AFE;
Xn_vect_imag = 256'h0507F41010080FFE03FE0C0BF0F90BFB09F0F9F60903F901FD0901F7FD05F306;
#100;

/*[(0.4375+0.25j), (0.125+0.375j), (-0.625+0.8125j), (0.5625+0.125j), (-0.3125-0.3125j), (-0.75-0.3125j), (-0.375+0.8125j), (0.6875+0.25j), (-0.625-0.25j), (0.8125-0.375j), (0.4375-0.6875j), (-0.0625-0.6875j), (-0.625+0.375j), (0.875+0.5625j), (-0.4375+0.125j), (-0.75-0.4375j), (0.5+0.6875j), (-0.9375+0.8125j), (0.1875+0.875j), (0.4375+0.1875j), (0.1875+0.8125j), (-0.375+0.5625j), -0.5j, (-0.1875-0.9375j), (-0.0625+0.1875j), (-0.0625-0.25j), (0.3125-0.3125j), (0.4375+0.5625j), (-0.0625-1j), (0.6875-0.0625j), (1-0.8125j), (-0.9375-0.9375j)]*/
Xn_vect_real = 256'h0702F609FBF4FA0BF60D07FFF60EF9F408F1030703FA00FDFFFF0507FF0B10F1;
Xn_vect_imag = 256'h04060D02FBFB0D04FCFAF5F5060902F90B0D0E030D09F8F103FCFB09F0FFF3F1;
#100;

/*[(0.875+0.75j), (-0.25-0.25j), (0.875-0.6875j), (-0.375-0.625j), (0.9375-0.0625j), (0.9375-0.25j), (-0.125+0.5j), (-0.1875-0.625j), (0.125-0.4375j), (0.875+0.1875j), (0.25+0.8125j), (-0.0625-0.8125j), (0.125+0.125j), (0.125+0.125j), (0.4375-0.875j), (-0.125+1j), 1j, 0.25j, (-0.125-0.5625j), (-0.9375+1j), (-0.4375-0.3125j), (-0.4375-0.5625j), (-0.1875-0.375j), (-0.5625-0.875j), (-0.75-0.4375j), (0.5625+0.4375j), (-0.6875+0.5j), (-0.5-1j), (0.0625+0.3125j), (-0.625-0.8125j), (-0.9375-0.8125j), (0.5625-1j)]*/
Xn_vect_real = 256'h0EFC0EFA0F0FFEFD020E04FF020207FE0000FEF1F9F9FDF7F409F5F801F6F109;
Xn_vect_imag = 256'h0CFCF5F6FFFC08F6F9030DF30202F2101004F710FBF7FAF2F90708F005F3F3F0;
#100;

/*[(0.9375-0.125j), (-0.8125+0j), (-0.1875-0.0625j), (-0.5625+0j), (0.0625-0.875j), (-0.8125-0.25j), (-0.6875+0.0625j), (0.625-0.6875j), (-0.125-0.5j), (-0.4375-0.9375j), (0.5625-0.8125j), (0.5625+1j), (-0.25-0.3125j), (-0.25-0.5625j), (0.125+0.9375j), (-0.125+0.25j), (-1-0.6875j), (-0.5+1j), (-0.4375-0.0625j), (-0.8125+0.8125j), (-0.1875-0.6875j), (-0.75+0.5625j), (-0.1875-1j), (0.5+0.3125j), (-0.6875+1j), (0.4375-0.875j), (-0.1875-0.625j), (0.3125+0.625j), (0.625+0.25j), (0.125+0.125j), (0.75-0.125j), 0.125j]*/
Xn_vect_real = 256'h0FF3FDF701F3F50AFEF90909FCFC02FEF0F8F9F3FDF4FD08F507FD050A020C00;
Xn_vect_imag = 256'hFE00FF00F2FC01F5F8F1F310FBF70F04F510FF0DF509F00510F2F60A0402FE02;
#100;

/*[(-0.75+0.625j), (0.25-0.375j), (-0.375+0.8125j), (0.1875-0.3125j), -0.25j, (-0.4375+0.6875j), (1-0.3125j), (-0.0625-0.125j), (-0.625+0.0625j), (-0.6875+0.9375j), (-0.75-1j), (0.75+0.4375j), (0.5625+0.1875j), (-0.875-0.25j), (-0.3125-0.75j), (-0.125-0.8125j), (0.75-0.4375j), (-0.4375-0.8125j), (-1+0.5j), (0.875-0.75j), (0.25+0j), (0.75+0.625j), (-0.4375+0.5625j), (0.5625+0.25j), (-1+0.4375j), (-0.5625+0.4375j), (-0.6875+0.875j), (-1-0.5j), (-0.5625+0.6875j), (0.6875-0.875j), (0.5625-0.6875j), (-0.1875+0.4375j)]*/
Xn_vect_real = 256'hF404FA0300F910FFF6F5F40C09F2FBFE0CF9F00E040CF909F0F7F5F0F70B09FD;
Xn_vect_imag = 256'h0AFA0DFBFC0BFBFE010FF00703FCF4F3F9F308F4000A090407070EF80BF2F507;
#100;

/*[(0.3125+0.6875j), (-0.8125-0.1875j), (-0.875-0.8125j), (0.4375+0j), (0.3125-0.375j), (0.3125-0.6875j), (-0.375-0.375j), (-0.0625-0.625j), -0.4375j, (0.3125+0.375j), (-0.5-0.875j), (-0.9375-0.6875j), (0.5625+0.3125j), (0.625+0j), (-0.25-1j), (-0.6875+0j), (0.875+0.9375j), (0.9375-0.5j), (0.875+0.1875j), (0.5625-0.0625j), (0.75+0.4375j), (0.8125-1j), (-0.6875+0.375j), (-0.1875-0.5625j), (1-0.1875j), (0.875-0.4375j), 0.5625j, (-0.5625-0.25j), (0.375+0.5625j), (0.9375+0.125j), (0.0625+0.875j), (0.8125-0.3125j)]*/
Xn_vect_real = 256'h05F3F2070505FAFF0005F8F1090AFCF50E0F0E090C0DF5FD100E00F7060F010D;
Xn_vect_imag = 256'h0BFDF300FAF5FAF6F906F2F50500F0000FF803FF07F006F7FDF909FC09020EFB;
#100;

/*[(0.125-0.3125j), (0.4375+0.125j), (-0.125+0.25j), (0.375+0.4375j), -0.75j, (-0.4375+0.125j), (-0.375-0.3125j), (0.9375+0.4375j), (0.125-1j), (-0.625+0.0625j), (0.5+0.75j), (0.25+0j), (-0.875-0.4375j), (0.5625-1j), (-0.8125-0.375j), (-0.625-0.5j), (-0.8125+0.625j), (-0.6875-0.0625j), (0.125+0.125j), (-0.8125+0.5625j), (-0.1875-0.625j), (-0.5+0.4375j), (0.3125+0.75j), (-0.1875-0.3125j), (0.25-0.3125j), (0.1875-0.125j), (0.875+0.0625j), (-0.4375+0.75j), (0.625+0.75j), (-0.0625+0.9375j), (-0.375-0.625j), (-0.1875+0.9375j)]*/
Xn_vect_real = 256'h0207FE0600F9FA0F02F60804F209F3F6F3F502F3FDF805FD04030EF90AFFFAFD;
Xn_vect_imag = 256'hFB020407F402FB07F0010C00F9F0FAF80AFF0209F6070CFBFBFE010C0C0FF60F;
#100;

/*[(-0.625-0.375j), (0.6875-0.5625j), (-0.6875-0.25j), (0.5625+0.25j), (0.625-0.0625j), (-0.6875-0.5j), (-0.6875+0.875j), (-0.25-0.1875j), (-0.875+0.875j), (-0.0625+0.625j), (-0.125+0.5j), (0.125-0.3125j), (-0.4375+0.125j), (0.4375+0.75j), (0.75-0.8125j), (0.0625-0.3125j), (-0.25+1j), (-0.8125+0.4375j), (0.25-0.5j), (0.375+0.75j), (0.6875-0.3125j), (0.375+0.75j), (-0.375+1j), (0.8125-0.4375j), (-0.875+0.5625j), (-0.375-0.375j), (-0.1875-1j), (-0.3125+0.375j), (0.125+0.3125j), (0.5625+0j), (0.375+0.5625j), (0.25-0.625j)]*/
Xn_vect_real = 256'hF60BF5090AF5F5FCF2FFFE02F9070C01FCF304060B06FA0DF2FAFDFB02090604;
Xn_vect_imag = 256'hFAF7FC04FFF80EFD0E0A08FB020CF3FB1007F80CFB0C10F909FAF006050009F6;
#100;

/*[(-0.5625+0j), (-0.9375-0.5625j), (-0.375+0.0625j), (0.375-0.75j), (0.375-0.3125j), (0.9375-0.9375j), (-0.3125+0.875j), (-0.5625+0.5625j), (0.5-0.3125j), (-0.4375+0.0625j), (-0.125-0.8125j), (-0.75-0.1875j), (0.8125+0.9375j), (-0.0625+0.5j), (0.25+0.25j), (-0.5625-0.5625j), (-0.1875-0.5625j), (0.1875+0.5j), (-0.5+0.9375j), (-0.25+0.1875j), (0.1875+0.375j), (0.25+0.1875j), (0.75-0.6875j), (0.1875+0.9375j), (0.9375-0.8125j), (-0.625-0.3125j), (1+0.5625j), (0.3125+0.375j), (0.5625-0.8125j), (-0.25+0.0625j), (0.5-0.6875j), (1+0.25j)]*/
Xn_vect_real = 256'hF7F1FA06060FFBF708F9FEF40DFF04F7FD03F8FC03040C030FF6100509FC0810;
Xn_vect_imag = 256'h00F701F4FBF10E09FB01F3FD0F0804F7F7080F030603F50FF3FB0906F301F504;
#100;

end

always @(Xn_vect_real,Xk_vect_imag)
$monitor("real=%h  imag=%h",Xk_vect_real,Xk_vect_imag);


//Expected output:
/*[-0.0625    -3.43750000e+00j -0.45419527-2.69144578e+00j
  1.71780271-7.01747321e+00j -2.99118476+6.92695451e+00j
 -1.80491748-4.71361156e+00j -3.99392064-1.56524327e-03j
  1.58086236+1.18583151e+00j  2.87137448-7.69978116e-01j
  5.25      -3.75000000e-01j  1.12675039-3.36455823e+00j
  2.64877829+1.90763544e+00j  4.92071909-1.31129009e+00j
  1.14590774-1.17287383e+00j  3.30738604-1.51259486e+00j
  2.43628062+1.43581377e+00j  2.87079922-4.08037527e+00j
  2.8125    -6.87500000e-01j -0.01978444-4.94642072e-01j
  3.20269242-5.42109218e-01j -5.14359669+2.28858632e+00j
 -2.07008252+4.21361156e+00j  4.36220483+4.15492083e+00j
  0.23607937-5.21508385e+00j -4.95435971+2.38952765e+00j
 -1.5       -5.00000000e+00j  4.46334584+3.20568524e-01j
  0.68072658-9.80530176e-02j  1.29464497+7.40040378e-01j
 -1.77090774-5.32712617e+00j  3.20821325+2.08931682e+00j
 -1.50322236+2.84343857e+00j  6.13160339-2.68346538e+00j]*/
//real=FFF91BD1E4C1192D54122A4E1234262D2D0033AEDF4503B1E8470A14E433E862  imag=C9D5906EB50012F4FACB1EECEEE816BFF5F9F8244342AD26B005FF0BAB212DD6
//real=fff71acee3c7172c5413294a1131262c2d0134b2df4305b8e8450d16e535ea60  imag=c9d29368b60310f5facd1ceeeceb17c0f5f8f520423db023b005000eac212ddc

/*[ 0.3125    +2.1875j      3.42998516+1.11144988j  3.98195044-0.53536385j
  2.77703413-2.00778865j -3.38756313-3.28553391j -0.40151311+0.68311284j
 -4.28857947+1.58765153j  0.49760017+3.91874088j -0.0625    -1.4375j
  0.98902814+4.49417423j  2.79309483+0.91988602j -7.21585561+0.07915634j
 -4.62760191-1.1061553j   2.84199027-5.10922175j -0.77619076-2.78615285j
 -2.01187708-8.20907281j  1.1875    +0.3125j      0.78081737-0.61724806j
  1.67705931+2.87115029j -2.43715375-3.706576j   -5.86243687+3.78553391j
 -2.87129137+2.14251984j -1.75951757+4.17275611j  3.39556331+3.94608185j
  0.0625    +3.9375j     -6.09627728-4.17771589j  6.04789542+4.24432754j
  0.1511015 -2.12519933j -1.62239809+2.6061553j  -1.17273918+0.97292889j
 -0.6757122 -3.47425479j -3.65641267+4.60465772j]*/
//real=05363F2CCAFABC07FF0F2C8DB62DF4E0130C1ADAA3D3E436019F6002E7EEF6C6  imag=2311F8E0CC0A193EE9470E01EFAFD48005F72DC53C22423F3FBE43DE290FC949


/*[ 0.5       +0.5j         1.78361831-2.51060324j  4.11370618+6.10212833j
  1.56387066+0.44285494j  1.41789322-2.30698052j  2.43551767+3.45342199j
  1.02676482+0.30050161j -0.42759236-3.06399661j  2.125     +0.25j
 -3.96973085-1.06756548j  7.05267995-3.42040557j  1.62119466-2.77090333j
  3.62392225+1.39016504j -1.79820226-0.416146j    1.04261242+1.61700584j
 -1.84823831-5.26876701j -0.625     +1.625j       0.83245954+2.35548397j
  6.24765294+0.16456088j  1.75278595+2.67793677j  2.83210678+4.05698052j
 -4.38043548+6.67908648j  5.54170109+3.44321682j  2.54223147-1.23392151j
 -4.25      +0.625j       0.23753647-2.34317925j -6.41403907-1.09628363j
 -2.90752119+5.72638325j -3.62392225+0.85983496j  0.8592366 -5.15049847j
 -5.61107832+0.88927573j  0.70326912-4.5095865j ]*/
//real=081C4119162610FA22C1701939E410E3F60D631C2DBA5828BC039AD2C70DA70B  imag=08D86107DC3704CF04EFCAD416FA19AC1A25022A406A37ED0ADBEF5B0DAE0EB8


/*[-0.5625    -4.37500000e+00j  3.3239718 -1.06505725e+01j
  0.82494016+8.09231021e-01j -0.26891048-5.58349342e+00j
  4.67883973+1.41107278e+00j -0.10531369+1.79779957e+00j
 -0.25201799+6.00902144e+00j  6.69386362+1.64796316e+00j
  3.5       -9.37500000e-01j  2.91609413+4.31608580e-01j
 -3.66725275+1.09318119e+01j -0.08524385+2.00901290e+00j
 -2.46024756+7.44257307e-01j  2.00575305+2.28077621e+00j
  5.77387188-7.92538693e-03j -0.42759065+5.62909019e+00j
  1.4375    +3.25000000e+00j  1.0586738 +3.63588744e+00j
  0.90361323-4.31595901e+00j  0.32559216-5.28417829e-01j
 -2.30383973-2.03607278e+00j -2.67433454-5.16944702e+00j
  2.40214425+4.10861925e+00j  0.23721659-1.72685202e+00j
 -0.625     +5.81250000e+00j  0.09034757-7.45350694e-01j
  4.68869936+1.82491606e+00j -0.00697173+1.29959749e+00j
 -1.66475244+3.13074269e+00j  0.38480789-5.80701633e-01j
  1.32600185+1.64028470e+00j  0.53204434+2.25309952e+00j]*/
//real=F7350DFC4AFFFC6B382EC6FFD9205CFA17100E05DCD62603F6014B00E6061508  imag=BA800CA7161C601AF1067F200B24005A343ABBF8E0AE41E55DF51D1432F71A24


/*[-3.37500000e+00-2.125j       1.95035276e-01-1.1990918j
 -2.47585861e+00+9.42165963j  2.56202194e+00+0.6624429j
  7.62081801e-04+0.14828644j -1.79861600e+00+0.77160775j
  3.10975577e+00-0.58000206j  4.37708908e+00+1.22078582j
 -3.75000000e+00+3.25j        1.13529816e+00+1.59042509j
  1.18842256e+00-9.08283235j -1.25951151e+00+4.92342161j
  2.24111652e-01+4.06770382j  3.82947785e-01-3.77971712j
  6.49960300e+00-0.85418361j  1.11121219e+00+3.31685986j
  1.62500000e+00-5.125j       4.30036689e+00+1.43184274j
  1.41780035e+00-2.8265433j   5.93427047e+00-0.29753927j
 -5.12576208e+00+2.97671356j  4.57439077e-01+1.82133117j
 -2.89134378e-01-3.48693968j  6.91947223e+00+1.50726902j
  3.00000000e+00-3.75j       -2.82004015e+00+1.00525109j
 -3.13036429e+00-0.76228398j  1.20991824e+00-0.08121846j
  4.00888348e-01-1.94270382j  1.64756897e+00-1.64164893j
 -3.20224397e-01-2.32887465j  6.64552737e+00-2.25202149j]*/
//real=CA03D92800E43146C41213EC030667111A44165EAE07FC6E30D3CE13061AFB6A  imag=DEED7F0A020CF7133419804E41C4F335AE16D3FC2F1DC918C410F4FFE1E6DBDC


/*[-3.6875    +0.3125j     -2.86591107+2.01398223j  3.61362442-7.54136019j
  3.97814343+4.4595354j  -1.66551452+4.96913104j -1.15664756+3.67387706j
  2.02589515+0.81431913j -9.43716645-2.17199267j  2.375     +3.625j
 -1.72534721-2.93817363j -3.3335597 -3.16308655j -1.03446968+1.22575686j
 -3.32192235-3.51830583j -5.29350775-2.1353379j   0.36040669+1.77868063j
  4.61275683+4.66605285j -3.0625    +2.3125j     -4.85959957-2.41391619j
  1.45223958+5.53247672j -4.40114961-3.22195294j  2.66551452+2.40586896j
  4.60213833+1.66007211j  8.24707562-1.11609583j -2.50640163+2.83037941j
 -1.125     -1.j         -4.05954979+4.32034064j  0.26769571+2.92197002j
 -1.27475719+0.10468017j -5.17807765-3.60669417j  0.35842462+1.31915568j
  0.36662254-1.72690393j  1.0630443 +3.60754092j]*/
//real=C5D3393FE6EE208026E5CBF0CBAC0549CFB317BA2A497FD8EEC004ECAE050511  imag=052088474F3A0DDE3AD1CE13C8DE1C4A25DA58CD261AEF2DF0452E01C715E539


/*[ 5.8125    -3.9375j     -5.44984446+4.99863976j -0.7365075 +1.98484333j
 -4.60751182+2.61354193j -0.40402913+0.77090774j  1.13367907+4.51242614j
 -4.10889891+2.67963028j -2.58916754+2.66867434j  6.125     -1.625j
  3.5129644 +0.34196392j  0.4852481 +6.67381097j  3.32022591+0.72871356j
  2.63518443+1.828966j    1.04076382+1.16458064j  0.17572673-0.81434997j
  2.84439504-0.083686j   -0.9375    +5.6875j     -6.8383367 +0.12742138j
  1.16588611+2.17676832j -2.87579302-0.89763498j -0.84597087-2.14590774j
 -1.40874187+1.69765073j  3.89919022+3.21941824j -1.62522364-6.53567777j
  5.75      +7.625j       0.75224598-3.35190854j -3.41462671-2.33542262j
  1.67564206-5.14652348j -0.63518443-0.203966j    0.75726976-3.49077403j
  4.03398196+4.41530145j  1.357433  -3.3474076j ]*/
//real=5DA9F5B7FA12BFD7623807352A10022DF19312D2F3EA3EE65C0CCA1AF60C4015  imag=C14F1F290C482A2AE6056A0B1D12F3FF5B0222F2DE1B33987ACBDBAEFDC946CB


/*[-2.4375    +1.375j       1.04311334+2.7088363j  -3.88991651+1.56349319j
 -2.62400596-0.87837977j  2.58210678-3.18121843j  2.04097891-4.51734765j
  0.96850165+1.44141326j  0.77784728+0.38978492j -2.6875    -2.25j
  2.80782828+1.76225257j -0.57411858-0.06489778j -3.03095399-2.72468837j
 -1.35983496+4.45526695j -4.57478575-3.45353732j -0.29733451+0.81355779j
  0.61829619-8.7939828j   1.1875    -4.25j       -0.31140264-0.05600726j
 -3.73140384-0.73659023j  3.33221849+2.70197273j  1.16789322-1.94378157j
 -1.81231777-3.147185j    5.23124581+4.93879056j  6.20161866+1.19145731j
  0.9375    -3.125j      -1.4788788 -0.94756719j -2.80456108+5.48799482j
  0.33746009-2.6417978j  -1.89016504+0.91973305j  4.28546444+1.15055555j
 -3.40241296-0.44376161j  7.38751925+2.25563378j]*/
//real=D910C2D729200F0CD52CF7D0EBB7FC0913FCC53512E453630FE9D405E244CA76  imag=162B19F2CEB81706DC1CFFD547C90D80BC00F52BE1CE4F13CEF157D60E12F924


/*[-0.5625    +3.125j       0.25204695-1.11899148j  4.21754587-2.60878594j
 -0.69508708+0.13353138j -6.05805826+1.30989809j -0.60298992-5.36180938j
 -0.89828764+1.94445597j -0.12769006-2.268903j    0.6875    +3.25j
 -1.60788183-3.69006624j -0.71886078-1.39356952j  3.60126048-4.85285897j
  1.282932  +4.63464556j -4.18181952-1.84023172j  1.20982877-2.45903531j
 -3.76758214+2.6755538j  -4.0625    +1.875j      -0.61411717+2.52293934j
  1.47592003-2.35460241j -4.7413741 +2.47598606j -6.94194174+4.31510191j
 -3.13697924-2.28909941j  4.0081226 +6.30967011j  3.76323584-1.61269074j
 -2.5625    +0.25j        3.31094232-0.2086778j  -4.72460512-3.39304213j
 -2.15223617-2.72632838j -2.782932  -2.25964556j  6.08079841+0.98593668j
  2.43033628-2.54509076j -1.38052677-4.82429015j]*/
//real=F70443F5A0F7F2FE0BE7F53914BE13C4BFF717B591CE403CD734B5DED46126EA  imag=32EFD70214AB1FDC34C5EAB34AE3D92A1E28DB2745DC64E704FDCAD5DC0FD8B3


/*[ 2.625     -0.6875j      0.93515225-0.42540494j -2.4001767 +0.27514485j
 -2.78616468-1.25951599j -3.07842712+2.49448052j -1.30748307+8.21593094j
  4.15099078+0.87614753j -1.98763684+5.72306124j  0.125     -1.3125j
 -4.31302131-0.12434859j -1.2189715 +1.86741769j  0.47139274+7.21278926j
 -1.80805826-1.91345148j -1.42652283-0.3800298j  -6.28802464-1.69458101j
 -5.1261644 -1.12474425j  5.        -1.3125j      1.86409664+1.39638662j
 -1.48110487+6.2755541j   2.77066123-3.92034671j  2.57842712-3.86948052j
 -0.05627947+3.22168262j -3.71640835+0.65678447j -1.69980824-3.06304641j
  2.75      -2.6875j      4.84219954-4.97836107j -3.89974694-2.91811663j
 -0.77390877+4.12392769j -2.69194174-4.21154852j  0.46185825+1.07414422j
 -2.64655779-0.83835099j  2.13162897-6.69212482j]*/
//real=2A0EDAD4CFEC42E102BBED07E4EA9CAE501DE92C2900C5E52C4DC2F4D507D622  imag=F5FA04EC277F0E5BEBFF1D73E2FAE5EFEB1664C2C3330ACFD5B1D241BD11F395


endmodule