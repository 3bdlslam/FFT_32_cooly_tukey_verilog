`timescale 1ns / 1ps

module complex_mul_test;
// Inputs
reg [3:-4] a;
reg [3:-4] aj;
reg [3:-4] b;
reg [3:-4] bj;

// Outputs
wire [3:-4] c;
wire [3:-4] cj;

// Instantiate the Unit Under Test (UUT)
complex_mul uut (
.a(a),
.aj(aj),
.b(b),
.bj(bj),
.c(c),
.cj(cj)
);
initial begin
// Initialize Inputs

//-1.0+j-0.375
a=0'hF0;
aj=0'hFA;
//0.8125+j-0.5
b=0'h0D;
bj=0'hF8;
#100;

//0.125+j-0.3125
a=0'h02;
aj=0'hFB;
//0.375+j-0.3125
b=0'h06;
bj=0'hFB;
#100;

//0.125+j-0.625
a=0'h02;
aj=0'hF6;
//-0.625+j0.8125
b=0'hF6;
bj=0'h0D;
#100;

//-0.25+j-0.25
a=0'hFC;
aj=0'hFC;
//0.1875+j-0.6875
b=0'h03;
bj=0'hF5;
#100;

//0.5+j0.75
a=0'h08;
aj=0'h0C;
//0.5625+j0.6875
b=0'h09;
bj=0'h0B;
#100;

//0.9375+j-0.1875
a=0'h0F;
aj=0'hFD;
//0.125+j-0.4375
b=0'h02;
bj=0'hF9;
#100;

//1.0+j0.125
a=0'h10;
aj=0'h02;
//0.6875+j0.25
b=0'h0B;
bj=0'h04;
#100;

//-0.75+j0.9375
a=0'hF4;
aj=0'h0F;
//0.6875+j0.75
b=0'h0B;
bj=0'h0C;
#100;

//0.75+j-0.875
a=0'h0C;
aj=0'hF2;
//0.75+j-1.0
b=0'h0C;
bj=0'hF0;
#100;

//0.5+j0.3125
a=0'h08;
aj=0'h05;
//-0.875+j0.25
b=0'hF2;
bj=0'h04;
#100;
end

always @(a,aj,b,bj)
$monitor("['%h','%h'],\n",c,cj);

/*Expected output:
[
(-1+0.1953125j)
['0'hF0','0'h03'],
(-0.05078125-0.15625j)
['0'h00','0'hFE'],
(0.4296875+0.4921875j)
['0'h06','0'h07'],
(-0.21875+0.125j)
['0'hFD','0'h02'],
(-0.234375+0.765625j)
['0'hFD','0'h0C'],
(0.03515625-0.43359375j)
['0'h00','0'hFA'],
(0.65625+0.3359375j)
['0'h0A','0'h05'],
(-1.21875+0.08203125j)
['0'hED','0'h01'],
(-0.3125-1.40625j)
['0'hFB','0'hEA'],
(-0.515625-0.1484375j)
['0'hF8','0'hFE'],
]*/

endmodule