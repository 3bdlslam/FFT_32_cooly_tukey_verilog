`timescale 1ns / 1ps

module Test_FFT;

// Inputs
reg [255:0] Xn_vect_real;
reg [255:0] Xn_vect_imag;
reg clk1,clk2,rst;
// Outputs
wire [255:0] Xk_vect_real;
wire [255:0] Xk_vect_imag;

// Instantiate the Unit Under Test (UUT)
FFT uut (
.Xn_vect_real(Xn_vect_real),
.Xn_vect_imag(Xn_vect_imag),
.Xk_vect_real(Xk_vect_real),
.Xk_vect_imag(Xk_vect_imag),
.clk1(clk1),.clk2(clk2),.rst(rst)
);

initial begin;
clk1<=0;
clk2<=1;
rst<=0;
#1 rst<=1;
#1 rst<=0;
end

always begin; #0.06172839506172839; clk1<=~clk1;
end
always begin; #5; clk2<=~clk2;
end

initial begin;

#10;
Xn_vect_real=  256'h00_00_00_00_00_FF_01_00_00_01_00_FF_01_00_00_00_00_01_00_01_00_01_FF_00_00_01_00_00_00_00_00_00;
Xn_vect_imag=  256'h00_00_00_00_00_00_FF_01_FF_00_01_00_00_01_00_00_00_00_01_00_00_00_00_01_FF_FF_FF_01_00_00_01_00;
#10;
Xn_vect_real=  256'hFF_00_00_00_FF_00_00_00_00_00_00_00_00_01_01_01_00_FF_00_01_01_00_00_00_01_00_00_01_00_00_FF_00;
Xn_vect_imag=  256'h00_01_00_00_00_00_01_00_00_00_00_00_01_00_FF_00_00_00_00_00_00_00_FF_00_00_01_00_FF_00_00_00_00;
#10;
Xn_vect_real=  256'h00_00_00_00_FF_00_01_00_01_00_01_00_00_00_00_01_00_00_00_00_00_00_FF_01_01_FF_01_01_00_FF_00_00;
Xn_vect_imag=  256'h00_01_00_00_00_00_FF_01_01_00_00_01_01_FF_01_01_FF_FF_01_FF_00_00_00_00_00_01_01_FF_00_00_00_00;
#10;
Xn_vect_real=  256'h01_00_FF_01_01_00_00_00_FF_00_FF_01_00_00_FF_00_00_FF_01_FF_01_00_01_00_FF_00_FF_00_01_00_00_00;
Xn_vect_imag=  256'h00_00_00_00_00_00_00_FF_00_00_00_01_01_FF_00_01_FF_00_00_FF_00_00_00_00_01_00_00_00_00_FF_01_01;
#10;
Xn_vect_real=  256'hFF_01_00_00_FF_01_01_00_FF_00_FF_00_01_01_00_00_00_01_FF_00_00_00_00_01_00_00_00_FF_00_FF_00_00;
Xn_vect_imag=  256'h00_00_00_00_00_00_00_00_00_00_00_00_00_01_01_00_01_00_00_00_00_00_FF_00_00_FF_FF_FF_01_FF_FF_00;
#10;
Xn_vect_real=  256'hFF_FF_00_01_FF_01_00_00_FF_01_00_00_00_FF_00_01_00_01_00_FF_00_FF_00_00_00_00_00_00_00_00_01_FF;
Xn_vect_imag=  256'h00_01_00_00_00_01_00_00_00_00_01_00_00_00_00_01_00_00_00_00_00_00_01_FF_FF_00_00_00_FF_00_00_00;
#10;
Xn_vect_real=  256'h00_FF_00_00_00_FF_00_01_00_00_00_00_FF_00_FF_00_00_00_01_00_FF_FF_00_01_00_FF_00_00_00_01_00_FF;
Xn_vect_imag=  256'h00_00_00_00_00_00_00_FF_00_00_FF_FF_01_00_01_FF_00_00_00_00_01_FF_00_FF_00_00_00_00_01_00_01_00;
#10;
Xn_vect_real=  256'hFF_00_00_01_01_00_FF_FF_00_01_00_01_01_00_00_00_00_FF_01_00_FF_FF_FF_01_00_00_FF_00_00_00_00_00;
Xn_vect_imag=  256'h00_00_00_00_FF_01_00_01_00_00_01_00_00_00_FF_FF_00_00_00_00_00_00_01_FF_01_00_01_00_FF_00_00_00;
#10;
Xn_vect_real=  256'h00_FF_00_01_01_00_00_FF_00_00_01_FF_FF_01_FF_00_00_00_00_FF_00_FF_01_00_01_00_FF_FF_00_00_00_00;
Xn_vect_imag=  256'h00_00_FF_FF_00_FF_01_FF_00_00_00_00_00_00_01_00_01_FF_01_00_00_00_00_00_00_00_00_00_00_00_00_00;
#10;
Xn_vect_real=  256'h00_00_00_00_FF_00_FF_00_00_FF_00_FF_00_00_01_FF_00_00_01_01_00_01_FF_00_FF_00_FF_01_00_01_01_00;
Xn_vect_imag=  256'h00_00_01_00_FF_00_01_FF_01_01_00_00_00_00_00_00_00_00_FF_00_00_00_00_01_FF_FF_00_00_01_00_00_00;
end

always @(posedge clk2)
$monitor("real=%h  imag=%h\n\n",Xk_vect_real,Xk_vect_imag);
endmodule

/*
Expected Output:

real=04FFFFFD000200FDFEFE0606FA000002FE0100FD00FFFE000400FB03020101FD  imag=02000204FCFE0004FA0102FAFD050205FCFA07000000FEFC0002FFFF000003FE


real=03FD00000000FF0303FFFD000102FFFBFDFFFDFE02FE01FDFDFFFC06FDFFFEF9  imag=010301FF01FF01F805000300FEFF0000FF01FEFEFD0100FEFF00FF080002FE00


real=0400FA0005030002FE02FD030000FF040200FBFE0504FEF40001020002FC00FD  imag=040000020100FEFC0409FA00FFFDFFFE02FC0302F904FD03FA00FF040302FC01


real=0002FF05FBFB0101010400020000040000FE03FFFC00050407010602FB000402  imag=0101FE030300000002FFFB01FBFB02FD0306F906FF05F701FEFE03FE00030200


real=00020001FF040200FFF600FFFBFF0002FA00FDFEFE0200FFFFFC000101FF00F9  imag=FEFB02FB0302FB0101020000FEFBFDFE020205FD02FD00FF070303FEFD0405FD


real=FE0200FB00FCFEFFFE01FF05FE060100FE000204FE0300FAFAFD02F900FBFEFB  imag=02FF0301000205FFFC0101FEFE02FBF9FE03000502FEFFFFFC0103FE00000000


real=FCFFFDFD01FCFC00010002000700020400010000FD030502FB02FDFC02FF0001  imag=FF020402FC04F80006FCFDFF010003FD09FFFE00FB0201FFFE000101FDFB0301


real=FF00010000F9FC0204FEFF01FDFB0402FDF901000000FEFF0004FAFEFC020000  imag=01FDFEFEFE0702FE00FC03FC0402FFFF01FCFD050400FF02FAFD01FE0505F905


real=FD00FD00FFFAFC04010103000304FAFF0503FF01FFFC05000100FEFA03010103  imag=FFFCFFFD02050303FD04020002F705FC07FFFDFF000100FD0101FFFE000203FD


real=FF0104FFFC06FF01FE00FBFA040306FAFDFF030002030001FE00FAFDFE0206FE  imag=0105000700FC0002FEFBFF0200FDFC0801FE03FF000402F9000101FF00FDFFFE


*/
