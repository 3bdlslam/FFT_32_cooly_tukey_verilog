`timescale 1ns / 1ps


module test_FFT_32;
// Inputs
reg [255:0] Xn_vect_real;
reg [255:0] Xn_vect_imag;
reg clk;
// Outputs
wire [255:0] Xk_vect_real;
wire [255:0] Xk_vect_imag;
// Instantiate the Unit Under Test (UUT)
FFT_32 uut (
.Xn_vect_real(Xn_vect_real),
.Xn_vect_imag(Xn_vect_imag),
.Xk_vect_real(Xk_vect_real),
.Xk_vect_imag(Xk_vect_imag),
.clk(clk)
);

initial begin

/*[(0.3125-0.1875j), (0.8125+0.3125j), (0.6875-0.375j), (-0.5-0.75j), (0.5625-0.3125j), (-1+1j), (-0.1875-0.6875j), (-0.6875-0.75j), (0.8125-0.875j), (-0.875-0.25j), (0.3125-0.875j), (-0.8125+0.5625j), (0.8125+0.125j), (-0.25+0.5j), (0.4375+0.1875j), (-0.4375+1j), (0.625+0.1875j), (0.0625-0.875j), (0.875+0.625j), (-0.5-0.25j), (-0.625-0.8125j), (-0.5625+1j), (0.75+0.5625j), (0.0625-0.75j), (-0.3125-0.1875j), (-0.375+0.5625j), (-0.5625-0.5j), (-0.0625-0.0625j), (-0.5625-0.4375j), (0.3125-0.4375j), (-0.8125+0.0625j), (0.5625+0j)]*/
Xn_vect_real <= 256'h050D0BF809F0FDF50DF205F30DFC07F90A010EF8F6F70C01FBFAF7FFF705F309;
Xn_vect_imag <= 256'hFD05FAF4FB10F5F4F2FCF2090208031003F20AFCF31009F4FD09F8FFF9F90100;
#100;

/*[(-0.3125+0.6875j), (0.125-0.9375j), (0.375-0.8125j), (0.75-0.625j), (0.4375+0.375j), (0.5-0.3125j), (-0.5-0.625j), (-0.25-0.5j), (0.375-0.3125j), (-0.25+0.6875j), (0.75-0.6875j), (0.25-0.0625j), (0.4375-0.6875j), (-0.6875-0.3125j), (0.5-0.75j), (0.625+0.8125j), (-0.375-0.125j), (-0.4375+0.8125j), (0.5+0.6875j), (0.125+0.875j), (0.375+1j), (0.0625-1j), (0.125-0.375j), (0.0625+0.375j), (0.375-0.9375j), (0.9375+0.125j), (-0.0625-0.3125j), (0.1875+0.25j), (-0.375-0.0625j), (-0.5625+0.5625j), (-0.0625-0.75j), (-0.5625+0.5625j)]*/
Xn_vect_real <= 256'hFB02060C0708F8FC06FC0C0407F5080AFAF9080206010201060FFF03FAF7FFF7;
Xn_vect_imag <= 256'h0BF1F3F606FBF6F8FB0BF5FFF5FBF40DFE0D0B0E10F0FA06F102FB04FF09F409;
#100;

/*[(0.875+0.9375j), (-0.0625-0.9375j), (0.125+1j), (-0.1875-0.875j), (0.6875-0.625j), 0.9375j, (1+0.375j), (0.6875-0.3125j), (0.8125+0.3125j), (0.5625-0.3125j), (-0.625-0.25j), (0.625-0.375j), (-0.125+0.875j), (0.25+0.0625j), (-0.4375-0.3125j), (0.1875-0.4375j), (-0.5625-0.3125j), (0.75-0.375j), (0.9375-0.8125j), (-0.4375+0.125j), (-0.625-0.625j), (-0.0625+0.6875j), (-0.875+0.3125j), (0.875+0.3125j), (-0.125+0j), (0.625+0.125j), (-0.125+0.5625j), (0.5+0.625j), (0.1875-0.4375j), (0.3125-0.25j), (-1-0.3125j), (-0.125-0.9375j)]*/
Xn_vect_real <= 256'h0EFF02FD0B00100B0D09F60AFE04F903F70C0FF9F6FFF20EFE0AFE080305F0FE;
Xn_vect_imag <= 256'h0FF110F2F60F06FB05FBFCFA0E01FBF9FBFAF302F60B05050002090AF9FCFBF1;
#100;

/*[(0.1875-0.5625j), (-0.375-0.125j), (0.5625+0.9375j), (0.1875+0.125j), (-0.8125+0.125j), (0.0625+0.3125j), (0.75+0.0625j), (-0.3125+0.5j), -0.1875j, (0.6875+0.25j), (-0.625+0.125j), (0.25+0.8125j), (0.375-0.0625j), (-0.3125+0.375j), (0.1875+0.5625j), (-0.4375-0.6875j), (-0.6875-0.3125j), (0.5+0.5625j), (-0.75-1j), (0.875+0.6875j), (-0.1875+0.1875j), (0.9375-0.4375j), (0.25-1j), (-0.75+0.125j), (-0.9375+0.6875j), (-0.4375-0.4375j), (-0.8125+0.3125j), (-1-0.3125j), (1+0.3125j), (-1+0.625j), (-0.8125+0.125j), (0.75-0.75j)]*/
Xn_vect_real <= 256'h03FA0903F3010CFB000BF60406FB03F9F508F40EFD0F04F4F1F9F3F010F0F30C;
Xn_vect_imag <= 256'hF7FE0F0202050108FD04020DFF0609F5FB09F00B03F9F0020BF905FB050A02F4;
#100;

/*[(0.375-0.3125j), (0.4375+0j), (0.125-0.9375j), (0.3125+0.25j), (-1+0.5625j), (-1-0.5j), (-1-0.875j), (0.0625+1j), (0.4375-0.875j), (-0.75-0.375j), (-0.9375+0.4375j), (-0.125-0.875j), (0.875-0.5j), (0.75-0.625j), (0.0625+0.5625j), (-0.6875-0.375j), (-0.4375-0.4375j), (0.8125-0.6875j), (0.1875+0.75j), (-0.125+0.1875j), (1-0.8125j), -0.875j, (0.1875+0.875j), (-0.375-0.9375j), (-0.0625-0.5625j), (-0.1875+0.0625j), (0.5625-0.875j), (-0.125+1j), (-0.25+0.6875j), (-0.3125+0j), (-0.3125-0.9375j), (0.8125+0.75j)]*/
Xn_vect_real <= 256'h06070205F0F0F00107F4F1FE0E0C01F5F90D03FE100003FAFFFD09FEFCFBFB0D;
Xn_vect_imag <= 256'hFB00F10409F8F210F2FA07F2F8F609FAF9F50C03F3F20EF1F701F2100B00F10C;
#100;

/*[(-0.9375+0.5j), (0.9375-0.1875j), (0.3125+0.875j), (-0.125+0.875j), (0.1875+1j), (1+0.875j), (0.625+0.5j), (-0.125-0.6875j), (0.4375-0.375j), (-1-0.5625j), (0.75-0.0625j), (-1-0.4375j), (-0.5625+0.5625j), (0.1875-1j), (-0.1875-0.9375j), (-0.0625+0.8125j), (1+0.4375j), (-0.4375-0.625j), (-0.0625+0.8125j), (-0.875-0.8125j), (-0.375-0.375j), (-0.125-0.75j), (0.8125+0.5j), (1+0.6875j), (0.4375+0.3125j), (0.75+0.75j), (0.75+0.8125j), (0.75+0.9375j), (0.25+0.875j), (-0.375-0.4375j), (-0.8125-1j), (0.9375+0.8125j)]*/
Xn_vect_real <= 256'hF10F05FE03100AFE07F00CF0F703FDFF10F9FFF2FAFE0D10070C0C0C04FAF30F;
Xn_vect_imag <= 256'h08FD0E0E100E08F5FAF7FFF909F0F10D07F60DF3FAF4080B050C0D0F0EF9F00D;
#100;

/*[(0.0625-0.375j), (-1-0.3125j), (0.125+0.5625j), (0.125+0.625j), (0.5625+0.25j), (-1-0.8125j), (0.5-0.5625j), (0.1875-0.6875j), (0.1875-0.9375j), (0.1875+0.8125j), (-0.9375+1j), (-0.625+0.6875j), (0.8125-0.0625j), (0.875-0.5j), (-0.625-0.625j), (-0.4375-0.375j), (0.125+0.625j), (0.0625-0.8125j), (0.9375+0.75j), (-0.5-0.875j), (0.5625+0.125j), (0.5+0.75j), (-0.875-0.75j), (-0.0625-0.25j), (0.875+0.25j), (-0.75+0.0625j), (-0.0625-0.1875j), (-1+0.75j), (-0.1875-0.3125j), (0.875-0.625j), (-0.125-0.25j), (0.4375-0.4375j)]*/
Xn_vect_real <= 256'h01F0020209F008030303F1F60D0EF6F902010FF80908F2FF0EF4FFF0FD0EFE07;
Xn_vect_imag <= 256'hFAFB090A04F3F7F5F10D100BFFF8F6FA0AF30CF2020CF4FC0401FD0CFBF6FCF9;
#100;

/*[(-0.4375+0.75j), (0.375-0.8125j), (-0.25+0.75j), (0.375-0.25j), (0.25-0.5j), (-0.125+0.75j), (-0.375+0.6875j), (0.875-0.875j), (1-0.8125j), (0.75+0.5j), (-0.25-0.8125j), (0.625-0.75j), (0.3125-0.9375j), (0.6875-0.8125j), (-0.5625+0.6875j), (-0.1875+0j), (0.0625+0.875j), (-0.5625+0.875j), (-0.6875+0.9375j), (-0.6875+0.375j), (-0.3125+0.0625j), (0.375-0.3125j), (-0.1875-0.0625j), (0.875+0.8125j), (-0.875+0.625j), (0.8125+0.875j), (-0.8125+0.125j), (0.4375-0.25j), (0.125+0.375j), (-0.1875+0.4375j), (-1+0.6875j), (0.3125-0.4375j)]*/
Xn_vect_real <= 256'hF906FC0604FEFA0E100CFC0A050BF7FD01F7F5F5FB06FD0EF20DF30702FDF005;
Xn_vect_imag <= 256'h0CF30CFCF80C0BF2F308F3F4F1F30B000E0E0F0601FBFF0D0A0E02FC06070BF9;
#100;

/*[(0.8125+0.375j), (0.9375+0.6875j), (0.125-0.5j), (0.9375+0.125j), (0.9375-0.4375j), (0.9375+0.4375j), (-0.625+0.625j), (-0.5+0.0625j), (-1-0.125j), (0.5625-0.625j), (0.5-0.1875j), (-0.9375-0.5625j), (-0.4375+0.9375j), (1-0.375j), (0.125+0.8125j), (-0.0625+0.5625j), (0.125-0.3125j), (0.3125+1j), (1+0.1875j), (-0.625+0.875j), (0.875+0.5j), (0.375+0.375j), (0.75+0.125j), (-0.5+1j), (-0.875+0.5j), (-0.3125-0.75j), (-0.75-0.375j), (0.875+0j), (1-0.3125j), (1+0.375j), (-1+0.875j), (-0.5625-0.9375j)]*/
Xn_vect_real <= 256'h0D0F020F0F0FF6F8F00908F1F91002FF020510F60E060CF8F2FBF40E1010F0F7;
Xn_vect_imag <= 256'h060BF802F9070A01FEF6FDF70FFA0D09FB10030E0806021008F4FA00FB060EF1;
#100;

/*[(-0.875-0.3125j), (0.375-0.75j), (0.4375+0.9375j), (-0.5625-0.5625j), (-0.3125-0.1875j), (-0.125-0.0625j), (0.3125+0.25j), (0.8125-0.75j), (0.5-0.9375j), (-0.3125-0.5625j), (-0.5-0.9375j), (0.1875-0.0625j), 0.6875j, (-0.125+0.5j), (0.375-0.75j), (0.3125+0.6875j), (-0.5+0.5625j), (-0.5625+0.75j), (0.6875-0.125j), (-1+0.75j), (0.75-0.875j), (-0.125+0.5j), (-0.0625-0.0625j), (-0.25-0.75j), (-0.9375-0.5j), (0.9375+0j), (0.4375+0.0625j), (0.9375-0.5j), (0.875-0.375j), (-0.5625-0.25j), (-0.3125-0.75j), (0.75-0.9375j)]*/
Xn_vect_real <= 256'hF20607F7FBFE050D08FBF80300FE0605F8F70BF00CFEFFFCF10F070F0EF7FB0C;
Xn_vect_imag <= 256'hFBF40FF7FDFF04F4F1F7F1FF0B08F40B090CFE0CF208FFF4F80001F8FAFCF4F1;
#100;

end

always @(Xn_vect_real,Xk_vect_imag)
$monitor("real=%h  imag=%h",Xk_vect_real,Xk_vect_imag);


//Expected output:
/*[-1.125     -2.6875j     -1.53760282-3.70465469j  3.47042143+2.12109932j
  5.81640831-1.16458104j  0.13258252-2.20840774j -1.81622198+0.8878117j
 -2.05595681-0.7510911j   2.49802734+3.25514726j  2.9375    -2.j
  5.23007297-0.95836783j -4.8775149 -3.83239675j  0.88713894-2.61040285j
 -0.90295138+3.31196113j  0.95641308+1.02455489j -3.13270314+5.01352673j
 -2.61073827+5.26710659j  7.375     -4.3125j     -6.9406459 -6.45379822j
 -1.21521761-0.43175949j -1.42286095-2.12628084j -0.13258252+0.70840774j
 -4.04313135-2.94233199j  5.0862869 -4.46642332j -3.14471768+3.83109424j
 -2.6875    -1.j          1.72304948-2.30780046j  1.12231108+7.64305692j
 -0.2451524 +1.83019692j  5.90295138-0.31196113j -1.57193348+2.4545866j
  5.10237305+3.20398769j  1.22189471-2.28228029j]*/
//real=EEE8375D02E3E0272F53B20EF20FCED77691EDEAFEC051CED51B11FD5EE75113  imag=D5C521EEDD0EF434E0F1C3D734105054BB99FADE0BD1B93DF0DC7A1DFC2733DC


/*[ 3.4375    -2.375j      -4.28059284-3.25471496j -1.17083093+1.31077494j
 -5.34734553-5.35872365j  0.96024756-2.76830583j -2.64399025+0.06111847j
 -3.99194439+3.46911902j -0.48725002+2.75589006j -2.75      +5.0625j
  3.46787302-2.19704239j -3.6531316 +3.65732517j -2.80422174+2.48516373j
 -1.25942235-3.39222808j  3.0035151 -0.01007679j -4.92717584-0.35619417j
 -2.23923473+3.07624709j  1.6875    -5.j         -1.84628323+0.28500752j
  5.90458814+2.22843862j  3.35191837+3.7023783j   0.16475244-2.85669417j
  2.42416913+3.51545028j -2.60272553+2.00943437j  0.13700632+2.10121172j
  1.375     +2.0625j     -0.24785121+5.94187609j  1.66937439-2.94653873j
  1.13543533-0.05369211j -3.11557765+3.76722808j  5.62316027+2.15838178j
 -2.72815425+5.12764078j  1.75369199-2.20847513j]*/
//real=37BCEEAB0FD6C1F9D437C6D4EC30B2DD1BE35E350226D70216FD1A12CF59D51C  imag=DACC14ABD400372C51DD3A27CA00FB31B004233BD3382021215FD1003C2252DD


/*[ 4.625     -1.25j        0.50387617-1.88080164j -2.47798895-4.66491691j
 -0.69234823+1.15109804j  1.62185922-2.7476213j   3.26638705+4.30651973j
  2.16944981-1.24856947j  1.68661722+1.02097389j  3.9375    -0.6875j
  4.81128637-3.40918611j -3.43292401+0.2409961j   2.66973141+1.68308765j
 -2.78867469+5.89406791j -4.11534462+2.67437759j  3.7741883 +6.88004583j
 -0.17337004+6.70874867j -4.375     +2.625j       6.4288619 +0.90486509j
  0.38592095-1.51598586j  0.98268773+4.95060116j  1.00314078+2.9976213j
  5.44325628+1.33273008j  1.7813754 -0.86646931j  1.72965508-3.45600194j
  0.3125    -0.1875j      3.56448023-0.90561506j -2.72500798+7.18990667j
  0.65604561+1.84909663j  3.66367469+0.85593209j -5.90280339-0.52288968j
 -2.47501351-3.51500705j  2.14098123+3.59239591j]*/
//real=4A08D9F51934221A3F4CCA2AD4BF3CFEBA66060F10571C1B0539D50A3AA2D922  imag=ECE2B612D544ED10F5CA031A5E2A6E6B2A0EE84F2F15F3C9FDF2731D0DF8C839


/*[-2.6875    +1.9375j      1.69248041-2.44522677j -0.02644965-4.25238418j
  4.46332805+1.24686148j -0.39200487-2.11948052j  0.94698363-2.81345997j
  2.87171372-5.49222293j  3.99760676-1.21835713j  0.8125    -0.4375j
 -1.27023066+1.67067055j  4.12132943+7.08000959j -2.71245291+5.4624109j
 -1.11167479-2.23039322j -6.3750987 +1.39330026j  0.92673877-3.3805814j
  4.92963668+3.23170706j -1.9375    -1.3125j      1.93993849+2.96803741j
 -2.50908426+3.77751045j  1.79843773-3.45443792j -1.98299513+4.24448052j
  3.72871414-4.3563533j  -4.59658746-7.66463132j  2.7390453 -5.5010605j
 -0.4375    +0.5625j     -3.59962512-2.52406381j  0.41420448-2.60513585j
  2.21325027+2.14681597j -3.76332521-3.64460678j  2.9368378 -3.39290436j
  2.29813496+1.53743565j -3.42885188+3.58606014j]*/
//real=D51B0047FA0F2D3F0DEC41D5EF9A0E4EE11FD81CE13BB72BF9C70623C42E24CA  imag=1FD9BC13DFD3A9EDF91A7157DD16CA33EB2F3CC943BB86A809D8D722C6CA1839


/*[-0.6875     -5.25j       -2.28833708 +4.8513712j
  2.92624827 +1.73876551j  2.15330766 -2.76749837j
  0.76332521 -3.21338835j  6.73287273 -2.63102551j
 -1.63741503 -2.94251233j -3.74156255+11.42886341j
 -1.9375     -1.25j       -0.65840286 +7.91344841j
 -1.94083828 +0.4953438j   3.88587138 -3.25198992j
  0.20266504 -2.45082521j -1.69035019 +1.93607714j
 -3.36806563 -0.03217515j -1.42307129 -8.23810344j
  0.3125     -1.25j       -2.38703358 -4.24700479j
 -2.02459784 +0.5326811j   3.85739523 +2.21582008j
 -1.88832521 -3.03661165j -0.6779545  -8.83383703j
  0.75353155 +3.06751233j  0.92429669 +5.16796536j
  6.0625     -1.25j       -0.97473116 -0.29509659j
 -2.46081215 +2.48320959j  3.97259057 +1.53069744j
 -0.32766504 +0.20082521j  5.94393664 -1.69393285j
  4.2519491  +0.15717515j -0.6288277  -1.08575456j]*/
//real=F5DC2E220C6BE6C5E1F6E13E03E5CBEA05DAE03DE2F60C0E61F1D93FFB5F44F6  imag=AC4D1BD4CDD6D17FEC7E07CCD91E0080ECBD0823D0803152ECFC271803E502EF


/*[ 4.0625    +4.6875j      0.52212755+8.0494105j  -1.45830109-2.14256995j
  1.45788303-9.50497444j  6.35929608+1.16811643j -2.9147079 -2.50874179j
  4.45333663+3.21313939j  0.80667721+2.43554499j -5.875     +1.j
 -1.81791142+0.4259566j  -6.57482938+0.46864558j -5.37004237+2.69687853j
 -4.01462617+1.31824269j  0.13727159-1.90162653j -5.3119705 +0.16269297j
 -6.49327897+0.20593367j  1.1875    +4.1875j     -4.45154636-4.93358776j
 -1.52653387-0.61523578j -3.34404577+3.98898791j  3.26570392-6.16811643j
 -5.03688488-0.48077315j  6.24165344+0.18590913j -3.78040774-1.36622104j
  2.375     +1.875j       2.14162135+2.18829821j  3.05966434+5.78916015j
  1.37232163-0.99675599j  0.13962617-1.06824269j -9.57996993-0.33893607j
 -5.38301957+0.93825851j  5.35089298+3.04060638j]*/
//real=4108E91765D2470CA2E397ABC002AC9913B9E8CB34B063C4262230150280AA55  imag=4B7FDE8012D833261006072B15E2020343B2F73F9EF902EB1E235CF1EFFB0F30


/*[-0.1875    -2.5j        -0.93669174-0.96830284j  0.59926211-2.38826334j
  2.12560559+3.99005748j  6.11059704+0.407932j    1.24191258-1.76830955j
 -7.92303546+0.72243834j -2.39626249+1.696554j    3.1875    -2.j
 -3.81402931+3.09883386j  0.33841635-0.47669066j  9.54816644-2.59434345j
 -1.63051948+5.61135912j -2.57417045-0.48146883j -2.74403073+7.62818934j
  0.47792335-2.0244321j   4.0625    +1.5j         0.80760886-1.58593498j
  1.62561162+1.141943j   -4.4194409 -3.80336179j  1.51440296-3.657932j
 -0.55313798+3.55090166j  2.37493842-2.62040912j  3.66721796-3.33454061j
  4.9375    +1.25j       -2.82465475-4.97657656j -3.06329009+3.473011j
  1.13475616-6.81722597j -7.99448052-4.11135912j -1.3468372 +0.63085723j
  1.79212777+0.01978143j -1.13796611-0.61270755j]*/
//real=FDF20922611382DA33C3057FE6D7D507410C1ABA18F8253A4FD3CF1281EB1CEE  imag=D8F1DA3F06E40B1BE031F9D759F97AE018E712C4C638D7CB14B13793BF0A00F7


/*[ 0.75      +3.5625j     -5.17486037-4.00186573j -1.96203132+3.83639509j
  1.02737919-6.43277836j  0.31954365+3.90349026j -4.24133322-4.62766895j
 -0.71701137-3.1335701j   3.16176672+4.82476145j  7.125     -2.0625j
 -0.96159955-2.27260031j -2.26072419+1.32640145j -4.88018956+4.55155306j
 -0.15533009+1.67861652j -2.58947159-2.40815069j  2.58709621+7.30630163j
 -1.55028484+4.07635564j -8.75      +3.3125j     -1.88544623-0.41563817j
  2.27269149+3.61703203j -1.15148894+3.2200817j  -3.56954365+0.72150974j
  0.89888572+2.55949205j  3.00254528-0.25183754j  1.97927783-1.51114852j
  1.375     -3.0625j     -3.97073453-1.3098958j   0.45006402+0.47017143j
  2.39033828+1.41850292j  0.90533009+3.44638348j  2.42455977-3.52367242j
 -7.37263011+1.32910601j  6.52320132+3.85267212j]*/
//real=0CAEE11005BDF53272F1DCB2FED729E880E224EEC70E301F16C107260E268B68  imag=39C03D9A3EB6CE4DDFDC15481ADA744135FA39330B28FCE8CFEC071637C8153D


/*[ 5.        +4.9375j     -0.40378117-2.74417691j  7.62225397-0.56433728j
 -1.10092729-0.4409577j  -9.76278634-2.09597087j -4.82845307-3.08470511j
  5.41685151-2.34963026j  9.63449494+0.79018862j  1.3125    -6.625j
  4.15165697+0.52880078j  6.1749879 -1.34877491j  2.22995192+2.70440128j
  2.07712617+1.50758252j  3.20741202+1.48158147j  6.36565479+1.7177863j
 -5.43312152-1.70289794j -1.875     +0.4375j     -1.91625369+2.34408429j
 -3.56419571-4.24004133j  3.45417348+4.9907039j  -3.48721366-1.65402913j
 -2.84145185+6.356922j   -0.16945342-0.81350556j  1.07079902-3.748024j
  1.3125    +5.75j        3.54490205+0.8231948j  -1.23304616-0.09684649j
 -2.69195533+5.07212416j -2.07712617+1.24241748j -0.41403127+0.79429867j
  1.88694712+5.19534951j  3.33658476-3.16553831j]*/
//real=50FA79EF80B3567F15426223213365AAE2E2C737C9D3FE111538EDD5DFFA1E35  imag=4FD5F7F9DFCFDB0C9608EB2B18171BE50725BD4FE665F3C55C0DFF51130C53CE


/*[ 1.5625    -5.3125j      0.97257967-4.37335508j -0.10046371+5.62352021j
  0.18987417-1.90100981j  0.64406791-2.55751939j  3.53600571-3.88935471j
  3.89048068+0.80321382j -1.91784308-2.43403368j  0.375     +1.125j
  2.89159184-1.5796014j  -9.16756003+3.2748945j  -1.26955486+1.84594952j
 -6.71729121+2.65479121j -3.89528448-3.22175168j  0.84576168+2.91348169j
 -4.60296961+5.50847368j  0.1875    -1.3125j     -1.57273316+5.63036826j
  1.66264805-3.31806386j  2.02188313+3.44548374j -4.39406791+0.18251939j
 -1.73856547-2.57228595j  0.34327654-0.24775747j -0.42659765-1.97460673j
 -4.125     -2.25j       -1.12202097-4.50799439j -1.6446243 +2.91964914j
  4.78787512+5.40031427j -2.03270879-2.02979121j -5.57157315-3.98602504j
 -3.32951889+1.53106195j  1.71733278-5.390571j  ]*/
//real=190FFF030A383EE2062E80EC95C20DB703E71A20BAE505FABEEFE64CE0A7CB1B  imag=ABBB59E2D8C20CDA12E7341D2ACD2E58EB5ACB3702D7FDE1DCB82E56E0C118AA


endmodule