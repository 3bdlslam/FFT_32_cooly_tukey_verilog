`timescale 1ns / 1ps

module complex_mul_test;
// Inputs
reg [3:-4] a;
reg [3:-4] aj;
reg [3:-4] b;
reg [3:-4] bj;

// Outputs
wire [3:-4] c;
wire [3:-4] cj;

// Instantiate the Unit Under Test (UUT)
complex_mul uut (
.a(a),
.aj(aj),
.b(b),
.bj(bj),
.c(c),
.cj(cj)
);
initial begin
// Initialize Inputs

//0.1875+j0.25
a=0'h03;
aj=0'h04;
//0.75+j-0.875
b=0'h0C;
bj=0'hF2;
#100;

//-0.375+j0.4375
a=0'hFA;
aj=0'h07;
//0.0625+j-0.125
b=0'h01;
bj=0'hFE;
#100;

//-1.0+j-1.0
a=0'hF0;
aj=0'hF0;
//-0.75+j-0.6875
b=0'hF4;
bj=0'hF5;
#100;

//-0.1875+j0.0
a=0'hFD;
aj=0'h00;
//0.875+j0.875
b=0'h0E;
bj=0'h0E;
#100;

//-0.5+j-0.625
a=0'hF8;
aj=0'hF6;
//0.625+j0.625
b=0'h0A;
bj=0'h0A;
#100;

//0.0625+j-0.625
a=0'h01;
aj=0'hF6;
//-0.75+j-0.5625
b=0'hF4;
bj=0'hF7;
#100;

//-0.1875+j0.875
a=0'hFD;
aj=0'h0E;
//1.0+j-0.625
b=0'h10;
bj=0'hF6;
#100;

//0.3125+j-0.5
a=0'h05;
aj=0'hF8;
//-0.8125+j0.0625
b=0'hF3;
bj=0'h01;
#100;

//0.3125+j0.75
a=0'h05;
aj=0'h0C;
//-1.0+j0.875
b=0'hF0;
bj=0'h0E;
#100;

//0.125+j-0.625
a=0'h02;
aj=0'hF6;
//0.4375+j-0.25
b=0'h07;
bj=0'hFC;
#100;
end

always @(a,aj,b,bj)
$monitor("['%h','%h'],\n",c,cj);

/*Expected output:
[
(0.359375+0.0234375j)
['0'h05','0'h00'],
(0.03125+0.07421875j)
['0'h00','0'h01'],
(0.0625+1.4375j)
['0'h01','0'h17'],
(-0.1640625-0.1640625j)
['0'hFE','0'hFE'],
(0.078125-0.703125j)
['0'h01','0'hF5'],
(-0.3984375+0.43359375j)
['0'hFA','0'h06'],
(0.359375+0.9921875j)
['0'h05','0'h0F'],
(-0.22265625+0.42578125j)
['0'hFD','0'h06'],
(-0.96875-0.4765625j)
['0'hF1','0'hF9'],
(-0.1015625-0.3046875j)
['0'hFF','0'hFC'],
]*/

endmodule