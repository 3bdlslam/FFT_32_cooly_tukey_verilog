`timescale 1ns / 1ps

module Test_FFT;

// Inputs
reg [255:0] Xn_vect_real;
reg [255:0] Xn_vect_imag;
reg clk1,clk2,rst;
// Outputs
wire [255:0] Xk_vect_real;
wire [255:0] Xk_vect_imag;

// Instantiate the Unit Under Test (UUT)
FFT uut (
.Xn_vect_real(Xn_vect_real),
.Xn_vect_imag(Xn_vect_imag),
.Xk_vect_real(Xk_vect_real),
.Xk_vect_imag(Xk_vect_imag),
.clk1(clk1),.clk2(clk2),.rst(rst)
);

initial begin;
clk1<=0;
clk2<=1;
rst<=0;
#1 rst<=1;
#1 rst<=0;
end

always begin; #0.06172839506172839; clk1<=~clk1;
end
always begin; #5; clk2<=~clk2;
end

initial begin;

#10;
Xn_vect_real=  256'hFF_00_FF_00_01_00_01_00_00_00_01_01_FF_00_01_00_01_FF_00_01_00_00_00_00_00_FF_01_FF_00_00_00_00;
Xn_vect_imag=  256'h00_00_01_01_FF_00_00_FF_01_01_01_01_01_00_01_00_00_00_FF_01_00_00_FF_01_FF_00_00_00_00_00_00_01;
#10;
Xn_vect_real=  256'hFF_00_01_00_00_00_FF_00_00_FF_01_00_FF_00_01_00_00_00_01_00_01_01_FF_01_00_00_FF_01_01_00_00_00;
Xn_vect_imag=  256'hFF_00_00_00_00_00_01_00_01_01_00_00_00_00_01_00_00_00_FF_FF_00_FF_00_FF_01_01_00_00_FF_00_00_00;
#10;
Xn_vect_real=  256'h00_00_01_00_01_01_FF_00_FF_00_00_00_00_00_00_01_00_FF_00_00_FF_00_01_01_00_00_00_01_00_01_FF_00;
Xn_vect_imag=  256'hFF_01_00_00_01_FF_00_00_00_00_00_01_00_00_00_00_00_00_FF_00_FF_00_01_FF_00_01_00_00_00_01_00_FF;
#10;
Xn_vect_real=  256'h00_FF_01_FF_00_00_00_00_00_01_00_00_00_00_00_00_00_00_FF_01_00_01_00_00_00_00_FF_00_FF_FF_00_00;
Xn_vect_imag=  256'h00_FF_01_00_00_00_FF_FF_00_00_00_00_00_01_01_00_00_00_FF_00_01_FF_00_FF_00_00_00_00_00_01_00_00;
#10;
Xn_vect_real=  256'hFF_00_00_00_00_00_00_00_00_00_01_00_00_00_00_01_00_00_00_00_01_00_00_01_00_00_FF_00_00_01_00_00;
Xn_vect_imag=  256'hFF_00_00_01_00_00_00_00_00_01_FF_FF_00_00_FF_00_00_00_00_00_00_01_00_00_01_FF_FF_00_00_00_00_00;
#10;
Xn_vect_real=  256'h00_01_01_FF_00_01_01_FF_00_00_FF_00_00_00_00_01_00_00_00_00_FF_FF_00_00_01_01_00_00_00_00_01_00;
Xn_vect_imag=  256'h00_00_00_00_01_01_00_FF_00_00_00_00_00_01_FF_00_00_00_00_00_00_00_01_00_00_00_00_00_00_00_01_FF;
#10;
Xn_vect_real=  256'hFF_00_00_FF_00_00_FF_00_00_00_00_00_00_00_00_FF_01_00_00_00_01_00_00_00_00_01_00_FF_FF_FF_00_00;
Xn_vect_imag=  256'h01_00_FF_01_00_00_01_00_01_00_FF_00_00_00_00_00_00_00_01_00_00_01_00_01_00_01_00_FF_00_00_00_01;
#10;
Xn_vect_real=  256'h00_FF_01_01_00_00_00_FF_00_00_01_FF_FF_00_00_00_00_00_00_01_00_FF_00_00_00_00_00_01_00_00_00_01;
Xn_vect_imag=  256'h00_00_00_00_00_01_00_00_00_01_01_00_00_FF_00_FF_FF_00_00_01_FF_00_00_00_01_FF_00_00_00_00_FF_01;
#10;
Xn_vect_real=  256'h00_00_00_01_00_00_00_00_00_00_00_00_00_01_FF_FF_FF_01_01_00_00_00_00_FF_00_00_00_00_00_00_00_00;
Xn_vect_imag=  256'hFF_00_00_01_01_FF_00_00_00_01_00_00_00_00_01_01_FF_FF_00_FF_00_01_00_01_00_00_00_00_01_FF_00_00;
#10;
Xn_vect_real=  256'h00_FF_01_FF_00_00_FF_FF_00_FF_00_00_00_00_01_00_01_FF_01_FF_00_00_00_00_01_00_00_00_00_00_00_01;
Xn_vect_imag=  256'h00_FF_00_00_FF_FF_FF_00_00_00_FF_00_00_FF_FF_00_00_00_00_00_FF_FF_00_FF_FF_00_00_00_00_00_FF_00;
end

always @(posedge clk2)
$monitor("real=%h  imag=%h\n\n",Xk_vect_real,Xk_vect_imag);
endmodule

/*
Expected Output:

real=0201FBFF0100FF01FA0000F803F801FA0404FAF701040502000003FDFBFE02F9  imag=06FD0006010002FD02FAFD0300FF00FFFC0101FE010203FEFC03FAFEFE040102


real=03020002FCFEFA010200FAFC04FE00FEFFFF0601FBFEFA02FC0001FDFEFE04FA  imag=0003FBFE02FEFEFA0103FB0204FEFD0002FAFE03FC0001FAFD00FE0305FDFDFD


real=0303FD0100FD020502040100050000FEFB000504FBFD00FCFC0300FAFDFC0201  imag=0002FEFA00FCFFFB010003FC04020001FE00FBFBFBFD0008FDFE00FEFE05FF00


real=FEFDFA050102FD0002FB00F801FF0006FE0306030103FEFEFEFF04FF010102FD  imag=FFFE0000FEFE0000010003000008000303FEFF000200FFFD0100FA00FC000601


real=03FD0400FDFD00FE01FCFD05FE000000FDFCFE03FDFC0301FF01FEFB0002FBFE  imag=FE00000101FCFDFB04FEFD0102FD0001FCFEFD00FF0100FD0204FCFCFE000000


real=030303FF0300FFFF0200FD000003FE04010100FDFFFEFCF9FA01000405FB0003  imag=020100FDFE0000FDFDFA04FE000101030203FE0204FEFD01030601FBFB03FF00


real=FCFA0201FF00FFFA01FEFCFBFF0303FC020001FAFEFD02FE010000040502FBFD  imag=0601FE0001040101FF03FF0700FC00FFFE0000FC0001030405FFFC0005010100


real=010503FC02FBFE05FCFB00FE01FD01000100FB0903FF04FFFE02FE00FD000000  imag=0004FC03FD000406030400020200FF01FEFCFCFF01FEFDFCFB05FD000301FD00


real=00010005FC06FBFFFC00FF030104FF00FE00FDFF00FD0104020100FDFFFC0100  imag=02FFFB02FAFFFC06FC05FE00FAFA01FF000300FEFA03FD0002FE00FA0200FF00


real=FFFF00FE050001FEFD02F7FC02FD01FE09FC0300020000FE0303FEFEFE020500  imag=F40304FC030002FF0202030205020300FE00FE00FBFF000000FFFFFE0001FFFD


*/
