`timescale 1ns / 1ps

module complex_mul_test;
// Inputs
reg [3:-4] a;
reg [3:-4] aj;
reg [3:-4] b;
reg [3:-4] bj;

// Outputs
wire [3:-4] c;
wire [3:-4] cj;

// Instantiate the Unit Under Test (UUT)
complex_mul uut (
.a(a),
.aj(aj),
.b(b),
.bj(bj),
.c(c),
.cj(cj)
);
initial begin
// Initialize Inputs

//2.5625+j-1.875
a=0'h29;
aj=0'hE2;
//1.0625+j-0.3125
b=0'h11;
bj=0'hFB;
#100;

//2.6875+j-5.0
a=0'h2B;
aj=0'hB0;
//0.3125+j0.9375
b=0'h05;
bj=0'h0F;
#100;

//-0.8125+j-0.4375
a=0'hF3;
aj=0'hF9;
//1.4375+j-3.5
b=0'h17;
bj=0'hC8;
#100;

//0.125+j-1.9375
a=0'h02;
aj=0'hE1;
//-3.4375+j-3.1875
b=0'hC9;
bj=0'hCD;
#100;

//-2.4375+j-4.6875
a=0'hD9;
aj=0'hB5;
//-1.625+j0.125
b=0'hE6;
bj=0'h02;
#100;

//0.875+j0.25
a=0'h0E;
aj=0'h04;
//-1.5625+j2.1875
b=0'hE7;
bj=0'h23;
#100;

//0.25+j-0.375
a=0'h04;
aj=0'hFA;
//-0.875+j-1.9375
b=0'hF2;
bj=0'hE1;
#100;

//1.375+j-0.375
a=0'h16;
aj=0'hFA;
//0.3125+j5.5
b=0'h05;
bj=0'h58;
#100;

//-1.0625+j0.0
a=0'hEF;
aj=0'h00;
//-1.375+j0.9375
b=0'hEA;
bj=0'h0F;
#100;

//-3.3125+j-0.1875
a=0'hCB;
aj=0'hFD;
//-1.4375+j2.4375
b=0'hE9;
bj=0'h27;
#100;

//-1.625+j3.6875
a=0'hE6;
aj=0'h3B;
//-0.75+j2.4375
b=0'hF4;
bj=0'h27;
#100;

//-1.25+j2.8125
a=0'hEC;
aj=0'h2D;
//0.5625+j1.0
b=0'h09;
bj=0'h10;
#100;

//1.1875+j1.0
a=0'h13;
aj=0'h10;
//-3.4375+j1.4375
b=0'hC9;
bj=0'h17;
#100;

//-2.9375+j7.1875
a=0'hD1;
aj=0'h73;
//0.375+j0.3125
b=0'h06;
bj=0'h05;
#100;

//-0.625+j1.75
a=0'hF6;
aj=0'h1C;
//3.25+j1.0
b=0'h34;
bj=0'h10;
#100;

//-0.125+j-0.0625
a=0'hFE;
aj=0'hFF;
//7.5625+j-1.0
b=0'h79;
bj=0'hF0;
#100;

//0.125+j2.875
a=0'h02;
aj=0'h2E;
//-0.0625+j0.8125
b=0'hFF;
bj=0'h0D;
#100;

//-1.625+j0.1875
a=0'hE6;
aj=0'h03;
//4.375+j4.25
b=0'h46;
bj=0'h44;
#100;

//-2.0+j0.3125
a=0'hE0;
aj=0'h05;
//2.1875+j0.5625
b=0'h23;
bj=0'h09;
#100;

//0.125+j-0.3125
a=0'h02;
aj=0'hFB;
//-2.5+j6.6875
b=0'hD8;
bj=0'h6B;
#100;

//1.5625+j-0.8125
a=0'h19;
aj=0'hF3;
//-2.875+j-3.8125
b=0'hD2;
bj=0'hC3;
#100;

//0.3125+j0.1875
a=0'h05;
aj=0'h03;
//3.8125+j3.625
b=0'h3D;
bj=0'h3A;
#100;

//-2.875+j-3.8125
a=0'hD2;
aj=0'hC3;
//0.6875+j0.0
b=0'h0B;
bj=0'h00;
#100;

//3.3125+j-0.625
a=0'h35;
aj=0'hF6;
//-1.8125+j-0.625
b=0'hE3;
bj=0'hF6;
#100;

//1.3125+j-0.875
a=0'h15;
aj=0'hF2;
//-0.5625+j2.75
b=0'hF7;
bj=0'h2C;
#100;

//3.9375+j-1.125
a=0'h3F;
aj=0'hEE;
//0.1875+j-0.6875
b=0'h03;
bj=0'hF5;
#100;
end

always @(a,aj,b,bj)
$monitor("['%h','%h'],\n",c,cj);

/*Expected output:
[
(2.13671875-2.79296875j)
['0'h22','0'hD4'],

(5.52734375+0.95703125j)
['0'h58','0'h0F'],

(-2.69921875+2.21484375j)
['0'hD5','0'h23'],

(-6.60546875+6.26171875j)
['0'h97','0'h64'],


(4.546875+7.3125j)
['0'h48','0'h75'],


(-1.9140625+1.5234375j)
['0'hE2','0'h18'],


(-0.9453125-0.15625j)
['0'hF1','0'hFE'],

(2.4921875+7.4453125j)
['0'h27','0'h77'],

(1.4609375-0.99609375j)
['0'h17','0'hF1'],


(5.21875-7.8046875j)
['0'h53','0'h84'],


(-7.76953125-6.7265625j)
['0'h84','0'h95'],


(-3.515625+0.33203125j)
['0'hC8','0'h05'],
(-5.51953125-1.73046875j)
['0'hA8','0'hE5'],
(-3.34765625+1.77734375j)
['0'hCB','0'h1C'],
(-3.78125+5.0625j)
['0'hC4','0'h51'],
(-1.0078125-0.34765625j)
['0'hF0','0'hFB'],
(-2.34375-0.078125j)
['0'hDB','0'hFF'],
(-7.90625-6.0859375j)
['0'h82','0'h9F'],
(-4.55078125-0.44140625j)
['0'hB8','0'hF9'],
(1.77734375+1.6171875j)
['0'h1C','0'h19'],
(-7.58984375-3.62109375j)
['0'h87','0'hC7'],
(0.51171875+1.84765625j)
['0'h08','0'h1D'],
(-1.9765625-2.62109375j)
['0'hE1','0'hD7'],
(-6.39453125-0.9375j)
['0'h9A','0'hF1'],
(1.66796875+4.1015625j)
['0'h1A','0'h41'],
(-0.03515625-2.91796875j)
['0'h00','0'hD2'],
]*/

endmodule